
`include "dump_file_agent.svh"
`include "csv_file_dump.svh"
`include "sample_agent.svh"
`include "loop_sample_agent.svh"
`include "sample_manager.svh"
`include "nodf_module_interface.svh"
`include "nodf_module_monitor.svh"
`include "pp_loop_interface.svh"
`include "pp_loop_monitor.svh"
`include "seq_loop_interface.svh"
`include "seq_loop_monitor.svh"
`include "upc_loop_interface.svh"
`include "upc_loop_monitor.svh"
`timescale 1ns/1ps

// top module for dataflow related monitors
module dataflow_monitor(
input logic clock,
input logic reset,
input logic finish
);



    nodf_module_intf module_intf_1(clock,reset);
    assign module_intf_1.ap_start = AESL_inst_TOP.ap_start;
    assign module_intf_1.ap_ready = AESL_inst_TOP.ap_ready;
    assign module_intf_1.ap_done = AESL_inst_TOP.ap_done;
    assign module_intf_1.ap_continue = 1'b1;
    assign module_intf_1.finish = finish;
    csv_file_dump mstatus_csv_dumper_1;
    nodf_module_monitor module_monitor_1;
    nodf_module_intf module_intf_2(clock,reset);
    assign module_intf_2.ap_start = AESL_inst_TOP.grp_TOP_Pipeline_VITIS_LOOP_461_1_fu_303.ap_start;
    assign module_intf_2.ap_ready = AESL_inst_TOP.grp_TOP_Pipeline_VITIS_LOOP_461_1_fu_303.ap_ready;
    assign module_intf_2.ap_done = AESL_inst_TOP.grp_TOP_Pipeline_VITIS_LOOP_461_1_fu_303.ap_done;
    assign module_intf_2.ap_continue = 1'b1;
    assign module_intf_2.finish = finish;
    csv_file_dump mstatus_csv_dumper_2;
    nodf_module_monitor module_monitor_2;
    nodf_module_intf module_intf_3(clock,reset);
    assign module_intf_3.ap_start = AESL_inst_TOP.grp_Rayleigh_fu_311.ap_start;
    assign module_intf_3.ap_ready = AESL_inst_TOP.grp_Rayleigh_fu_311.ap_ready;
    assign module_intf_3.ap_done = AESL_inst_TOP.grp_Rayleigh_fu_311.ap_done;
    assign module_intf_3.ap_continue = 1'b1;
    assign module_intf_3.finish = finish;
    csv_file_dump mstatus_csv_dumper_3;
    nodf_module_monitor module_monitor_3;
    nodf_module_intf module_intf_4(clock,reset);
    assign module_intf_4.ap_start = AESL_inst_TOP.grp_Rayleigh_fu_311.grp_seedInitialization_fu_40.ap_start;
    assign module_intf_4.ap_ready = AESL_inst_TOP.grp_Rayleigh_fu_311.grp_seedInitialization_fu_40.ap_ready;
    assign module_intf_4.ap_done = AESL_inst_TOP.grp_Rayleigh_fu_311.grp_seedInitialization_fu_40.ap_done;
    assign module_intf_4.ap_continue = 1'b1;
    assign module_intf_4.finish = finish;
    csv_file_dump mstatus_csv_dumper_4;
    nodf_module_monitor module_monitor_4;
    nodf_module_intf module_intf_5(clock,reset);
    assign module_intf_5.ap_start = AESL_inst_TOP.grp_Rayleigh_fu_311.grp_seedInitialization_fu_40.grp_seedInitialization_Pipeline_SEED_INIT_LOOP_fu_94.ap_start;
    assign module_intf_5.ap_ready = AESL_inst_TOP.grp_Rayleigh_fu_311.grp_seedInitialization_fu_40.grp_seedInitialization_Pipeline_SEED_INIT_LOOP_fu_94.ap_ready;
    assign module_intf_5.ap_done = AESL_inst_TOP.grp_Rayleigh_fu_311.grp_seedInitialization_fu_40.grp_seedInitialization_Pipeline_SEED_INIT_LOOP_fu_94.ap_done;
    assign module_intf_5.ap_continue = 1'b1;
    assign module_intf_5.finish = finish;
    csv_file_dump mstatus_csv_dumper_5;
    nodf_module_monitor module_monitor_5;
    nodf_module_intf module_intf_6(clock,reset);
    assign module_intf_6.ap_start = AESL_inst_TOP.grp_Rayleigh_fu_311.grp_Rayleigh_Pipeline_VITIS_LOOP_28_1_VITIS_LOOP_29_2_fu_54.ap_start;
    assign module_intf_6.ap_ready = AESL_inst_TOP.grp_Rayleigh_fu_311.grp_Rayleigh_Pipeline_VITIS_LOOP_28_1_VITIS_LOOP_29_2_fu_54.ap_ready;
    assign module_intf_6.ap_done = AESL_inst_TOP.grp_Rayleigh_fu_311.grp_Rayleigh_Pipeline_VITIS_LOOP_28_1_VITIS_LOOP_29_2_fu_54.ap_done;
    assign module_intf_6.ap_continue = 1'b1;
    assign module_intf_6.finish = finish;
    csv_file_dump mstatus_csv_dumper_6;
    nodf_module_monitor module_monitor_6;
    nodf_module_intf module_intf_7(clock,reset);
    assign module_intf_7.ap_start = AESL_inst_TOP.grp_Rayleigh_fu_311.grp_Rayleigh_Pipeline_VITIS_LOOP_40_3_VITIS_LOOP_41_4_fu_66.ap_start;
    assign module_intf_7.ap_ready = AESL_inst_TOP.grp_Rayleigh_fu_311.grp_Rayleigh_Pipeline_VITIS_LOOP_40_3_VITIS_LOOP_41_4_fu_66.ap_ready;
    assign module_intf_7.ap_done = AESL_inst_TOP.grp_Rayleigh_fu_311.grp_Rayleigh_Pipeline_VITIS_LOOP_40_3_VITIS_LOOP_41_4_fu_66.ap_done;
    assign module_intf_7.ap_continue = 1'b1;
    assign module_intf_7.finish = finish;
    csv_file_dump mstatus_csv_dumper_7;
    nodf_module_monitor module_monitor_7;
    nodf_module_intf module_intf_8(clock,reset);
    assign module_intf_8.ap_start = AESL_inst_TOP.grp_Rayleigh_fu_311.grp_Rayleigh_Pipeline_VITIS_LOOP_69_6_fu_74.ap_start;
    assign module_intf_8.ap_ready = AESL_inst_TOP.grp_Rayleigh_fu_311.grp_Rayleigh_Pipeline_VITIS_LOOP_69_6_fu_74.ap_ready;
    assign module_intf_8.ap_done = AESL_inst_TOP.grp_Rayleigh_fu_311.grp_Rayleigh_Pipeline_VITIS_LOOP_69_6_fu_74.ap_done;
    assign module_intf_8.ap_continue = 1'b1;
    assign module_intf_8.finish = finish;
    csv_file_dump mstatus_csv_dumper_8;
    nodf_module_monitor module_monitor_8;
    nodf_module_intf module_intf_9(clock,reset);
    assign module_intf_9.ap_start = AESL_inst_TOP.grp_AWGN_fu_319.ap_start;
    assign module_intf_9.ap_ready = AESL_inst_TOP.grp_AWGN_fu_319.ap_ready;
    assign module_intf_9.ap_done = AESL_inst_TOP.grp_AWGN_fu_319.ap_done;
    assign module_intf_9.ap_continue = 1'b1;
    assign module_intf_9.finish = finish;
    csv_file_dump mstatus_csv_dumper_9;
    nodf_module_monitor module_monitor_9;
    nodf_module_intf module_intf_10(clock,reset);
    assign module_intf_10.ap_start = AESL_inst_TOP.grp_AWGN_fu_319.grp_seedInitialization_fu_432.ap_start;
    assign module_intf_10.ap_ready = AESL_inst_TOP.grp_AWGN_fu_319.grp_seedInitialization_fu_432.ap_ready;
    assign module_intf_10.ap_done = AESL_inst_TOP.grp_AWGN_fu_319.grp_seedInitialization_fu_432.ap_done;
    assign module_intf_10.ap_continue = 1'b1;
    assign module_intf_10.finish = finish;
    csv_file_dump mstatus_csv_dumper_10;
    nodf_module_monitor module_monitor_10;
    nodf_module_intf module_intf_11(clock,reset);
    assign module_intf_11.ap_start = AESL_inst_TOP.grp_AWGN_fu_319.grp_seedInitialization_fu_432.grp_seedInitialization_Pipeline_SEED_INIT_LOOP_fu_94.ap_start;
    assign module_intf_11.ap_ready = AESL_inst_TOP.grp_AWGN_fu_319.grp_seedInitialization_fu_432.grp_seedInitialization_Pipeline_SEED_INIT_LOOP_fu_94.ap_ready;
    assign module_intf_11.ap_done = AESL_inst_TOP.grp_AWGN_fu_319.grp_seedInitialization_fu_432.grp_seedInitialization_Pipeline_SEED_INIT_LOOP_fu_94.ap_done;
    assign module_intf_11.ap_continue = 1'b1;
    assign module_intf_11.finish = finish;
    csv_file_dump mstatus_csv_dumper_11;
    nodf_module_monitor module_monitor_11;
    nodf_module_intf module_intf_12(clock,reset);
    assign module_intf_12.ap_start = AESL_inst_TOP.grp_TOP_Pipeline_VITIS_LOOP_482_2_VITIS_LOOP_483_3_fu_325.ap_start;
    assign module_intf_12.ap_ready = AESL_inst_TOP.grp_TOP_Pipeline_VITIS_LOOP_482_2_VITIS_LOOP_483_3_fu_325.ap_ready;
    assign module_intf_12.ap_done = AESL_inst_TOP.grp_TOP_Pipeline_VITIS_LOOP_482_2_VITIS_LOOP_483_3_fu_325.ap_done;
    assign module_intf_12.ap_continue = 1'b1;
    assign module_intf_12.finish = finish;
    csv_file_dump mstatus_csv_dumper_12;
    nodf_module_monitor module_monitor_12;
    nodf_module_intf module_intf_13(clock,reset);
    assign module_intf_13.ap_start = AESL_inst_TOP.grp_TOP_Pipeline_VITIS_LOOP_488_4_fu_346.ap_start;
    assign module_intf_13.ap_ready = AESL_inst_TOP.grp_TOP_Pipeline_VITIS_LOOP_488_4_fu_346.ap_ready;
    assign module_intf_13.ap_done = AESL_inst_TOP.grp_TOP_Pipeline_VITIS_LOOP_488_4_fu_346.ap_done;
    assign module_intf_13.ap_continue = 1'b1;
    assign module_intf_13.finish = finish;
    csv_file_dump mstatus_csv_dumper_13;
    nodf_module_monitor module_monitor_13;
    nodf_module_intf module_intf_14(clock,reset);
    assign module_intf_14.ap_start = AESL_inst_TOP.grp_TOP_Pipeline_VITIS_LOOP_492_5_VITIS_LOOP_493_6_fu_352.ap_start;
    assign module_intf_14.ap_ready = AESL_inst_TOP.grp_TOP_Pipeline_VITIS_LOOP_492_5_VITIS_LOOP_493_6_fu_352.ap_ready;
    assign module_intf_14.ap_done = AESL_inst_TOP.grp_TOP_Pipeline_VITIS_LOOP_492_5_VITIS_LOOP_493_6_fu_352.ap_done;
    assign module_intf_14.ap_continue = 1'b1;
    assign module_intf_14.finish = finish;
    csv_file_dump mstatus_csv_dumper_14;
    nodf_module_monitor module_monitor_14;
    nodf_module_intf module_intf_15(clock,reset);
    assign module_intf_15.ap_start = AESL_inst_TOP.grp_QRD_fu_389.ap_start;
    assign module_intf_15.ap_ready = AESL_inst_TOP.grp_QRD_fu_389.ap_ready;
    assign module_intf_15.ap_done = AESL_inst_TOP.grp_QRD_fu_389.ap_done;
    assign module_intf_15.ap_continue = 1'b1;
    assign module_intf_15.finish = finish;
    csv_file_dump mstatus_csv_dumper_15;
    nodf_module_monitor module_monitor_15;
    nodf_module_intf module_intf_16(clock,reset);
    assign module_intf_16.ap_start = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_V_fu_3293.ap_start;
    assign module_intf_16.ap_ready = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_V_fu_3293.ap_ready;
    assign module_intf_16.ap_done = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_V_fu_3293.ap_done;
    assign module_intf_16.ap_continue = 1'b1;
    assign module_intf_16.finish = finish;
    csv_file_dump mstatus_csv_dumper_16;
    nodf_module_monitor module_monitor_16;
    nodf_module_intf module_intf_17(clock,reset);
    assign module_intf_17.ap_start = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_V_fu_3293.grp_CORDIC_V_Pipeline_VITIS_LOOP_94_2_fu_173.ap_start;
    assign module_intf_17.ap_ready = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_V_fu_3293.grp_CORDIC_V_Pipeline_VITIS_LOOP_94_2_fu_173.ap_ready;
    assign module_intf_17.ap_done = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_V_fu_3293.grp_CORDIC_V_Pipeline_VITIS_LOOP_94_2_fu_173.ap_done;
    assign module_intf_17.ap_continue = 1'b1;
    assign module_intf_17.finish = finish;
    csv_file_dump mstatus_csv_dumper_17;
    nodf_module_monitor module_monitor_17;
    nodf_module_intf module_intf_18(clock,reset);
    assign module_intf_18.ap_start = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3308.ap_start;
    assign module_intf_18.ap_ready = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3308.ap_ready;
    assign module_intf_18.ap_done = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3308.ap_done;
    assign module_intf_18.ap_continue = 1'b1;
    assign module_intf_18.finish = finish;
    csv_file_dump mstatus_csv_dumper_18;
    nodf_module_monitor module_monitor_18;
    nodf_module_intf module_intf_19(clock,reset);
    assign module_intf_19.ap_start = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3308.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_start;
    assign module_intf_19.ap_ready = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3308.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_ready;
    assign module_intf_19.ap_done = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3308.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_done;
    assign module_intf_19.ap_continue = 1'b1;
    assign module_intf_19.finish = finish;
    csv_file_dump mstatus_csv_dumper_19;
    nodf_module_monitor module_monitor_19;
    nodf_module_intf module_intf_20(clock,reset);
    assign module_intf_20.ap_start = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3326.ap_start;
    assign module_intf_20.ap_ready = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3326.ap_ready;
    assign module_intf_20.ap_done = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3326.ap_done;
    assign module_intf_20.ap_continue = 1'b1;
    assign module_intf_20.finish = finish;
    csv_file_dump mstatus_csv_dumper_20;
    nodf_module_monitor module_monitor_20;
    nodf_module_intf module_intf_21(clock,reset);
    assign module_intf_21.ap_start = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3326.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_start;
    assign module_intf_21.ap_ready = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3326.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_ready;
    assign module_intf_21.ap_done = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3326.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_done;
    assign module_intf_21.ap_continue = 1'b1;
    assign module_intf_21.finish = finish;
    csv_file_dump mstatus_csv_dumper_21;
    nodf_module_monitor module_monitor_21;
    nodf_module_intf module_intf_22(clock,reset);
    assign module_intf_22.ap_start = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3335.ap_start;
    assign module_intf_22.ap_ready = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3335.ap_ready;
    assign module_intf_22.ap_done = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3335.ap_done;
    assign module_intf_22.ap_continue = 1'b1;
    assign module_intf_22.finish = finish;
    csv_file_dump mstatus_csv_dumper_22;
    nodf_module_monitor module_monitor_22;
    nodf_module_intf module_intf_23(clock,reset);
    assign module_intf_23.ap_start = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3335.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_start;
    assign module_intf_23.ap_ready = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3335.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_ready;
    assign module_intf_23.ap_done = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3335.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_done;
    assign module_intf_23.ap_continue = 1'b1;
    assign module_intf_23.finish = finish;
    csv_file_dump mstatus_csv_dumper_23;
    nodf_module_monitor module_monitor_23;
    nodf_module_intf module_intf_24(clock,reset);
    assign module_intf_24.ap_start = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3344.ap_start;
    assign module_intf_24.ap_ready = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3344.ap_ready;
    assign module_intf_24.ap_done = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3344.ap_done;
    assign module_intf_24.ap_continue = 1'b1;
    assign module_intf_24.finish = finish;
    csv_file_dump mstatus_csv_dumper_24;
    nodf_module_monitor module_monitor_24;
    nodf_module_intf module_intf_25(clock,reset);
    assign module_intf_25.ap_start = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3344.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_start;
    assign module_intf_25.ap_ready = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3344.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_ready;
    assign module_intf_25.ap_done = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3344.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_done;
    assign module_intf_25.ap_continue = 1'b1;
    assign module_intf_25.finish = finish;
    csv_file_dump mstatus_csv_dumper_25;
    nodf_module_monitor module_monitor_25;
    nodf_module_intf module_intf_26(clock,reset);
    assign module_intf_26.ap_start = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3353.ap_start;
    assign module_intf_26.ap_ready = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3353.ap_ready;
    assign module_intf_26.ap_done = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3353.ap_done;
    assign module_intf_26.ap_continue = 1'b1;
    assign module_intf_26.finish = finish;
    csv_file_dump mstatus_csv_dumper_26;
    nodf_module_monitor module_monitor_26;
    nodf_module_intf module_intf_27(clock,reset);
    assign module_intf_27.ap_start = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3353.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_start;
    assign module_intf_27.ap_ready = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3353.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_ready;
    assign module_intf_27.ap_done = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3353.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_done;
    assign module_intf_27.ap_continue = 1'b1;
    assign module_intf_27.finish = finish;
    csv_file_dump mstatus_csv_dumper_27;
    nodf_module_monitor module_monitor_27;
    nodf_module_intf module_intf_28(clock,reset);
    assign module_intf_28.ap_start = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3362.ap_start;
    assign module_intf_28.ap_ready = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3362.ap_ready;
    assign module_intf_28.ap_done = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3362.ap_done;
    assign module_intf_28.ap_continue = 1'b1;
    assign module_intf_28.finish = finish;
    csv_file_dump mstatus_csv_dumper_28;
    nodf_module_monitor module_monitor_28;
    nodf_module_intf module_intf_29(clock,reset);
    assign module_intf_29.ap_start = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3362.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_start;
    assign module_intf_29.ap_ready = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3362.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_ready;
    assign module_intf_29.ap_done = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3362.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_done;
    assign module_intf_29.ap_continue = 1'b1;
    assign module_intf_29.finish = finish;
    csv_file_dump mstatus_csv_dumper_29;
    nodf_module_monitor module_monitor_29;
    nodf_module_intf module_intf_30(clock,reset);
    assign module_intf_30.ap_start = AESL_inst_TOP.grp_QRD_fu_389.grp_QRD_Pipeline_LOOP_01_fu_3374.ap_start;
    assign module_intf_30.ap_ready = AESL_inst_TOP.grp_QRD_fu_389.grp_QRD_Pipeline_LOOP_01_fu_3374.ap_ready;
    assign module_intf_30.ap_done = AESL_inst_TOP.grp_QRD_fu_389.grp_QRD_Pipeline_LOOP_01_fu_3374.ap_done;
    assign module_intf_30.ap_continue = 1'b1;
    assign module_intf_30.finish = finish;
    csv_file_dump mstatus_csv_dumper_30;
    nodf_module_monitor module_monitor_30;
    nodf_module_intf module_intf_31(clock,reset);
    assign module_intf_31.ap_start = AESL_inst_TOP.grp_QRD_fu_389.grp_QRD_Pipeline_LOOP_02_VITIS_LOOP_251_6_fu_3469.ap_start;
    assign module_intf_31.ap_ready = AESL_inst_TOP.grp_QRD_fu_389.grp_QRD_Pipeline_LOOP_02_VITIS_LOOP_251_6_fu_3469.ap_ready;
    assign module_intf_31.ap_done = AESL_inst_TOP.grp_QRD_fu_389.grp_QRD_Pipeline_LOOP_02_VITIS_LOOP_251_6_fu_3469.ap_done;
    assign module_intf_31.ap_continue = 1'b1;
    assign module_intf_31.finish = finish;
    csv_file_dump mstatus_csv_dumper_31;
    nodf_module_monitor module_monitor_31;
    nodf_module_intf module_intf_32(clock,reset);
    assign module_intf_32.ap_start = AESL_inst_TOP.grp_QRD_fu_389.grp_QRD_Pipeline_VITIS_LOOP_268_8_fu_3539.ap_start;
    assign module_intf_32.ap_ready = AESL_inst_TOP.grp_QRD_fu_389.grp_QRD_Pipeline_VITIS_LOOP_268_8_fu_3539.ap_ready;
    assign module_intf_32.ap_done = AESL_inst_TOP.grp_QRD_fu_389.grp_QRD_Pipeline_VITIS_LOOP_268_8_fu_3539.ap_done;
    assign module_intf_32.ap_continue = 1'b1;
    assign module_intf_32.finish = finish;
    csv_file_dump mstatus_csv_dumper_32;
    nodf_module_monitor module_monitor_32;
    nodf_module_intf module_intf_33(clock,reset);
    assign module_intf_33.ap_start = AESL_inst_TOP.grp_QRD_fu_389.grp_QRD_Pipeline_VITIS_LOOP_316_9_VITIS_LOOP_317_10_fu_3674.ap_start;
    assign module_intf_33.ap_ready = AESL_inst_TOP.grp_QRD_fu_389.grp_QRD_Pipeline_VITIS_LOOP_316_9_VITIS_LOOP_317_10_fu_3674.ap_ready;
    assign module_intf_33.ap_done = AESL_inst_TOP.grp_QRD_fu_389.grp_QRD_Pipeline_VITIS_LOOP_316_9_VITIS_LOOP_317_10_fu_3674.ap_done;
    assign module_intf_33.ap_continue = 1'b1;
    assign module_intf_33.finish = finish;
    csv_file_dump mstatus_csv_dumper_33;
    nodf_module_monitor module_monitor_33;
    nodf_module_intf module_intf_34(clock,reset);
    assign module_intf_34.ap_start = AESL_inst_TOP.grp_TOP_Pipeline_VITIS_LOOP_433_1_fu_445.ap_start;
    assign module_intf_34.ap_ready = AESL_inst_TOP.grp_TOP_Pipeline_VITIS_LOOP_433_1_fu_445.ap_ready;
    assign module_intf_34.ap_done = AESL_inst_TOP.grp_TOP_Pipeline_VITIS_LOOP_433_1_fu_445.ap_done;
    assign module_intf_34.ap_continue = 1'b1;
    assign module_intf_34.finish = finish;
    csv_file_dump mstatus_csv_dumper_34;
    nodf_module_monitor module_monitor_34;
    nodf_module_intf module_intf_35(clock,reset);
    assign module_intf_35.ap_start = AESL_inst_TOP.grp_KBEST_fu_461.ap_start;
    assign module_intf_35.ap_ready = AESL_inst_TOP.grp_KBEST_fu_461.ap_ready;
    assign module_intf_35.ap_done = AESL_inst_TOP.grp_KBEST_fu_461.ap_done;
    assign module_intf_35.ap_continue = 1'b1;
    assign module_intf_35.finish = finish;
    csv_file_dump mstatus_csv_dumper_35;
    nodf_module_monitor module_monitor_35;
    nodf_module_intf module_intf_36(clock,reset);
    assign module_intf_36.ap_start = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_1_fu_903.ap_start;
    assign module_intf_36.ap_ready = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_1_fu_903.ap_ready;
    assign module_intf_36.ap_done = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_1_fu_903.ap_done;
    assign module_intf_36.ap_continue = 1'b1;
    assign module_intf_36.finish = finish;
    csv_file_dump mstatus_csv_dumper_36;
    nodf_module_monitor module_monitor_36;
    nodf_module_intf module_intf_37(clock,reset);
    assign module_intf_37.ap_start = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_VITIS_LOOP_347_1_fu_939.ap_start;
    assign module_intf_37.ap_ready = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_VITIS_LOOP_347_1_fu_939.ap_ready;
    assign module_intf_37.ap_done = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_VITIS_LOOP_347_1_fu_939.ap_done;
    assign module_intf_37.ap_continue = 1'b1;
    assign module_intf_37.finish = finish;
    csv_file_dump mstatus_csv_dumper_37;
    nodf_module_monitor module_monitor_37;
    nodf_module_intf module_intf_38(clock,reset);
    assign module_intf_38.ap_start = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_VITIS_LOOP_364_3_fu_947.ap_start;
    assign module_intf_38.ap_ready = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_VITIS_LOOP_364_3_fu_947.ap_ready;
    assign module_intf_38.ap_done = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_VITIS_LOOP_364_3_fu_947.ap_done;
    assign module_intf_38.ap_continue = 1'b1;
    assign module_intf_38.finish = finish;
    csv_file_dump mstatus_csv_dumper_38;
    nodf_module_monitor module_monitor_38;
    nodf_module_intf module_intf_39(clock,reset);
    assign module_intf_39.ap_start = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_VITIS_LOOP_420_10_fu_1009.ap_start;
    assign module_intf_39.ap_ready = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_VITIS_LOOP_420_10_fu_1009.ap_ready;
    assign module_intf_39.ap_done = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_VITIS_LOOP_420_10_fu_1009.ap_done;
    assign module_intf_39.ap_continue = 1'b1;
    assign module_intf_39.finish = finish;
    csv_file_dump mstatus_csv_dumper_39;
    nodf_module_monitor module_monitor_39;
    nodf_module_intf module_intf_40(clock,reset);
    assign module_intf_40.ap_start = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_VITIS_LOOP_373_5_fu_1016.ap_start;
    assign module_intf_40.ap_ready = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_VITIS_LOOP_373_5_fu_1016.ap_ready;
    assign module_intf_40.ap_done = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_VITIS_LOOP_373_5_fu_1016.ap_done;
    assign module_intf_40.ap_continue = 1'b1;
    assign module_intf_40.finish = finish;
    csv_file_dump mstatus_csv_dumper_40;
    nodf_module_monitor module_monitor_40;
    nodf_module_intf module_intf_41(clock,reset);
    assign module_intf_41.ap_start = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_VITIS_LOOP_391_6_VITIS_LOOP_392_7_fu_1058.ap_start;
    assign module_intf_41.ap_ready = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_VITIS_LOOP_391_6_VITIS_LOOP_392_7_fu_1058.ap_ready;
    assign module_intf_41.ap_done = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_VITIS_LOOP_391_6_VITIS_LOOP_392_7_fu_1058.ap_done;
    assign module_intf_41.ap_continue = 1'b1;
    assign module_intf_41.finish = finish;
    csv_file_dump mstatus_csv_dumper_41;
    nodf_module_monitor module_monitor_41;
    nodf_module_intf module_intf_42(clock,reset);
    assign module_intf_42.ap_start = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_VITIS_LOOP_410_9_fu_1136.ap_start;
    assign module_intf_42.ap_ready = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_VITIS_LOOP_410_9_fu_1136.ap_ready;
    assign module_intf_42.ap_done = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_VITIS_LOOP_410_9_fu_1136.ap_done;
    assign module_intf_42.ap_continue = 1'b1;
    assign module_intf_42.finish = finish;
    csv_file_dump mstatus_csv_dumper_42;
    nodf_module_monitor module_monitor_42;

    pp_loop_intf #(4) pp_loop_intf_1(clock,reset);
    assign pp_loop_intf_1.pre_loop_state0 = AESL_inst_TOP.grp_AWGN_fu_319.ap_ST_fsm_state2;
    assign pp_loop_intf_1.pre_states_valid = 1'b1;
    assign pp_loop_intf_1.post_loop_state0 = AESL_inst_TOP.grp_AWGN_fu_319.ap_ST_fsm_state33;
    assign pp_loop_intf_1.post_states_valid = 1'b1;
    assign pp_loop_intf_1.iter_start_state = AESL_inst_TOP.grp_AWGN_fu_319.ap_ST_fsm_pp0_stage0;
    assign pp_loop_intf_1.iter_start_enable = AESL_inst_TOP.grp_AWGN_fu_319.ap_enable_reg_pp0_iter0;
    assign pp_loop_intf_1.iter_start_block = AESL_inst_TOP.grp_AWGN_fu_319.ap_block_pp0_stage0_subdone;
    assign pp_loop_intf_1.iter_end_state = AESL_inst_TOP.grp_AWGN_fu_319.ap_ST_fsm_pp0_stage0;
    assign pp_loop_intf_1.iter_end_enable = AESL_inst_TOP.grp_AWGN_fu_319.ap_enable_reg_pp0_iter29;
    assign pp_loop_intf_1.iter_end_block = AESL_inst_TOP.grp_AWGN_fu_319.ap_block_pp0_stage0_subdone;
    assign pp_loop_intf_1.loop_quit_state = AESL_inst_TOP.grp_AWGN_fu_319.ap_ST_fsm_pp0_stage0;
    assign pp_loop_intf_1.quit_at_end = 1'b1;
    assign pp_loop_intf_1.cur_state = AESL_inst_TOP.grp_AWGN_fu_319.ap_CS_fsm;
    assign pp_loop_intf_1.finish = finish;
    csv_file_dump pp_loop_csv_dumper_1;
    pp_loop_monitor #(4) pp_loop_monitor_1;
    seq_loop_intf#(59) seq_loop_intf_1(clock,reset);
    assign seq_loop_intf_1.pre_loop_state0 = AESL_inst_TOP.grp_QRD_fu_389.ap_ST_fsm_state1;
    assign seq_loop_intf_1.pre_states_valid = 1'b1;
    assign seq_loop_intf_1.post_loop_state0 = AESL_inst_TOP.grp_QRD_fu_389.ap_ST_fsm_state12;
    assign seq_loop_intf_1.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_1.post_loop_state1 = 59'h0;
    assign seq_loop_intf_1.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_1.quit_loop_state0 = AESL_inst_TOP.grp_QRD_fu_389.ap_ST_fsm_state2;
    assign seq_loop_intf_1.quit_states_valid = 1'b1;
    assign seq_loop_intf_1.cur_state = AESL_inst_TOP.grp_QRD_fu_389.ap_CS_fsm;
    assign seq_loop_intf_1.iter_start_state = AESL_inst_TOP.grp_QRD_fu_389.ap_ST_fsm_state2;
    assign seq_loop_intf_1.iter_end_state0 = AESL_inst_TOP.grp_QRD_fu_389.ap_ST_fsm_state11;
    assign seq_loop_intf_1.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_1.one_state_loop = 1'b0;
    assign seq_loop_intf_1.one_state_block = 1'b0;
    assign seq_loop_intf_1.finish = finish;
    csv_file_dump seq_loop_csv_dumper_1;
    seq_loop_monitor #(59) seq_loop_monitor_1;
    seq_loop_intf#(59) seq_loop_intf_2(clock,reset);
    assign seq_loop_intf_2.pre_loop_state0 = AESL_inst_TOP.grp_QRD_fu_389.ap_ST_fsm_state2;
    assign seq_loop_intf_2.pre_states_valid = 1'b1;
    assign seq_loop_intf_2.post_loop_state0 = AESL_inst_TOP.grp_QRD_fu_389.ap_ST_fsm_state28;
    assign seq_loop_intf_2.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_2.post_loop_state1 = 59'h0;
    assign seq_loop_intf_2.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_2.quit_loop_state0 = AESL_inst_TOP.grp_QRD_fu_389.ap_ST_fsm_state12;
    assign seq_loop_intf_2.quit_states_valid = 1'b1;
    assign seq_loop_intf_2.cur_state = AESL_inst_TOP.grp_QRD_fu_389.ap_CS_fsm;
    assign seq_loop_intf_2.iter_start_state = AESL_inst_TOP.grp_QRD_fu_389.ap_ST_fsm_state12;
    assign seq_loop_intf_2.iter_end_state0 = AESL_inst_TOP.grp_QRD_fu_389.ap_ST_fsm_state27;
    assign seq_loop_intf_2.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_2.one_state_loop = 1'b0;
    assign seq_loop_intf_2.one_state_block = 1'b0;
    assign seq_loop_intf_2.finish = finish;
    csv_file_dump seq_loop_csv_dumper_2;
    seq_loop_monitor #(59) seq_loop_monitor_2;
    seq_loop_intf#(59) seq_loop_intf_3(clock,reset);
    assign seq_loop_intf_3.pre_loop_state0 = AESL_inst_TOP.grp_QRD_fu_389.ap_ST_fsm_state29;
    assign seq_loop_intf_3.pre_states_valid = 1'b1;
    assign seq_loop_intf_3.post_loop_state0 = AESL_inst_TOP.grp_QRD_fu_389.ap_ST_fsm_state38;
    assign seq_loop_intf_3.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_3.post_loop_state1 = 59'h0;
    assign seq_loop_intf_3.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_3.quit_loop_state0 = AESL_inst_TOP.grp_QRD_fu_389.ap_ST_fsm_state30;
    assign seq_loop_intf_3.quit_states_valid = 1'b1;
    assign seq_loop_intf_3.cur_state = AESL_inst_TOP.grp_QRD_fu_389.ap_CS_fsm;
    assign seq_loop_intf_3.iter_start_state = AESL_inst_TOP.grp_QRD_fu_389.ap_ST_fsm_state30;
    assign seq_loop_intf_3.iter_end_state0 = AESL_inst_TOP.grp_QRD_fu_389.ap_ST_fsm_state37;
    assign seq_loop_intf_3.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_3.one_state_loop = 1'b0;
    assign seq_loop_intf_3.one_state_block = 1'b0;
    assign seq_loop_intf_3.finish = finish;
    csv_file_dump seq_loop_csv_dumper_3;
    seq_loop_monitor #(59) seq_loop_monitor_3;
    seq_loop_intf#(59) seq_loop_intf_4(clock,reset);
    assign seq_loop_intf_4.pre_loop_state0 = AESL_inst_TOP.grp_QRD_fu_389.ap_ST_fsm_state40;
    assign seq_loop_intf_4.pre_states_valid = 1'b1;
    assign seq_loop_intf_4.post_loop_state0 = AESL_inst_TOP.grp_QRD_fu_389.ap_ST_fsm_state47;
    assign seq_loop_intf_4.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_4.post_loop_state1 = 59'h0;
    assign seq_loop_intf_4.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_4.quit_loop_state0 = AESL_inst_TOP.grp_QRD_fu_389.ap_ST_fsm_state41;
    assign seq_loop_intf_4.quit_states_valid = 1'b1;
    assign seq_loop_intf_4.cur_state = AESL_inst_TOP.grp_QRD_fu_389.ap_CS_fsm;
    assign seq_loop_intf_4.iter_start_state = AESL_inst_TOP.grp_QRD_fu_389.ap_ST_fsm_state41;
    assign seq_loop_intf_4.iter_end_state0 = AESL_inst_TOP.grp_QRD_fu_389.ap_ST_fsm_state46;
    assign seq_loop_intf_4.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_4.one_state_loop = 1'b0;
    assign seq_loop_intf_4.one_state_block = 1'b0;
    assign seq_loop_intf_4.finish = finish;
    csv_file_dump seq_loop_csv_dumper_4;
    seq_loop_monitor #(59) seq_loop_monitor_4;
    seq_loop_intf#(59) seq_loop_intf_5(clock,reset);
    assign seq_loop_intf_5.pre_loop_state0 = AESL_inst_TOP.grp_QRD_fu_389.ap_ST_fsm_state52;
    assign seq_loop_intf_5.pre_states_valid = 1'b1;
    assign seq_loop_intf_5.post_loop_state0 = AESL_inst_TOP.grp_QRD_fu_389.ap_ST_fsm_state55;
    assign seq_loop_intf_5.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_5.post_loop_state1 = 59'h0;
    assign seq_loop_intf_5.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_5.quit_loop_state0 = AESL_inst_TOP.grp_QRD_fu_389.ap_ST_fsm_state53;
    assign seq_loop_intf_5.quit_states_valid = 1'b1;
    assign seq_loop_intf_5.cur_state = AESL_inst_TOP.grp_QRD_fu_389.ap_CS_fsm;
    assign seq_loop_intf_5.iter_start_state = AESL_inst_TOP.grp_QRD_fu_389.ap_ST_fsm_state53;
    assign seq_loop_intf_5.iter_end_state0 = AESL_inst_TOP.grp_QRD_fu_389.ap_ST_fsm_state54;
    assign seq_loop_intf_5.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_5.one_state_loop = 1'b0;
    assign seq_loop_intf_5.one_state_block = 1'b0;
    assign seq_loop_intf_5.finish = finish;
    csv_file_dump seq_loop_csv_dumper_5;
    seq_loop_monitor #(59) seq_loop_monitor_5;
    seq_loop_intf#(7) seq_loop_intf_6(clock,reset);
    assign seq_loop_intf_6.pre_loop_state0 = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_V_fu_3293.ap_ST_fsm_state1;
    assign seq_loop_intf_6.pre_states_valid = 1'b1;
    assign seq_loop_intf_6.post_loop_state0 = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_V_fu_3293.ap_ST_fsm_state5;
    assign seq_loop_intf_6.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_6.post_loop_state1 = 7'h0;
    assign seq_loop_intf_6.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_6.quit_loop_state0 = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_V_fu_3293.ap_ST_fsm_state2;
    assign seq_loop_intf_6.quit_states_valid = 1'b1;
    assign seq_loop_intf_6.cur_state = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_V_fu_3293.ap_CS_fsm;
    assign seq_loop_intf_6.iter_start_state = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_V_fu_3293.ap_ST_fsm_state2;
    assign seq_loop_intf_6.iter_end_state0 = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_V_fu_3293.ap_ST_fsm_state4;
    assign seq_loop_intf_6.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_6.one_state_loop = 1'b0;
    assign seq_loop_intf_6.one_state_block = 1'b0;
    assign seq_loop_intf_6.finish = finish;
    csv_file_dump seq_loop_csv_dumper_6;
    seq_loop_monitor #(7) seq_loop_monitor_6;
    seq_loop_intf#(7) seq_loop_intf_7(clock,reset);
    assign seq_loop_intf_7.pre_loop_state0 = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3308.ap_ST_fsm_state1;
    assign seq_loop_intf_7.pre_states_valid = 1'b1;
    assign seq_loop_intf_7.post_loop_state0 = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3308.ap_ST_fsm_state5;
    assign seq_loop_intf_7.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_7.post_loop_state1 = 7'h0;
    assign seq_loop_intf_7.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_7.quit_loop_state0 = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3308.ap_ST_fsm_state2;
    assign seq_loop_intf_7.quit_states_valid = 1'b1;
    assign seq_loop_intf_7.cur_state = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3308.ap_CS_fsm;
    assign seq_loop_intf_7.iter_start_state = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3308.ap_ST_fsm_state2;
    assign seq_loop_intf_7.iter_end_state0 = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3308.ap_ST_fsm_state4;
    assign seq_loop_intf_7.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_7.one_state_loop = 1'b0;
    assign seq_loop_intf_7.one_state_block = 1'b0;
    assign seq_loop_intf_7.finish = finish;
    csv_file_dump seq_loop_csv_dumper_7;
    seq_loop_monitor #(7) seq_loop_monitor_7;
    seq_loop_intf#(7) seq_loop_intf_8(clock,reset);
    assign seq_loop_intf_8.pre_loop_state0 = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3326.ap_ST_fsm_state1;
    assign seq_loop_intf_8.pre_states_valid = 1'b1;
    assign seq_loop_intf_8.post_loop_state0 = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3326.ap_ST_fsm_state5;
    assign seq_loop_intf_8.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_8.post_loop_state1 = 7'h0;
    assign seq_loop_intf_8.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_8.quit_loop_state0 = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3326.ap_ST_fsm_state2;
    assign seq_loop_intf_8.quit_states_valid = 1'b1;
    assign seq_loop_intf_8.cur_state = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3326.ap_CS_fsm;
    assign seq_loop_intf_8.iter_start_state = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3326.ap_ST_fsm_state2;
    assign seq_loop_intf_8.iter_end_state0 = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3326.ap_ST_fsm_state4;
    assign seq_loop_intf_8.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_8.one_state_loop = 1'b0;
    assign seq_loop_intf_8.one_state_block = 1'b0;
    assign seq_loop_intf_8.finish = finish;
    csv_file_dump seq_loop_csv_dumper_8;
    seq_loop_monitor #(7) seq_loop_monitor_8;
    seq_loop_intf#(7) seq_loop_intf_9(clock,reset);
    assign seq_loop_intf_9.pre_loop_state0 = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3335.ap_ST_fsm_state1;
    assign seq_loop_intf_9.pre_states_valid = 1'b1;
    assign seq_loop_intf_9.post_loop_state0 = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3335.ap_ST_fsm_state5;
    assign seq_loop_intf_9.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_9.post_loop_state1 = 7'h0;
    assign seq_loop_intf_9.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_9.quit_loop_state0 = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3335.ap_ST_fsm_state2;
    assign seq_loop_intf_9.quit_states_valid = 1'b1;
    assign seq_loop_intf_9.cur_state = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3335.ap_CS_fsm;
    assign seq_loop_intf_9.iter_start_state = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3335.ap_ST_fsm_state2;
    assign seq_loop_intf_9.iter_end_state0 = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3335.ap_ST_fsm_state4;
    assign seq_loop_intf_9.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_9.one_state_loop = 1'b0;
    assign seq_loop_intf_9.one_state_block = 1'b0;
    assign seq_loop_intf_9.finish = finish;
    csv_file_dump seq_loop_csv_dumper_9;
    seq_loop_monitor #(7) seq_loop_monitor_9;
    seq_loop_intf#(7) seq_loop_intf_10(clock,reset);
    assign seq_loop_intf_10.pre_loop_state0 = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3344.ap_ST_fsm_state1;
    assign seq_loop_intf_10.pre_states_valid = 1'b1;
    assign seq_loop_intf_10.post_loop_state0 = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3344.ap_ST_fsm_state5;
    assign seq_loop_intf_10.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_10.post_loop_state1 = 7'h0;
    assign seq_loop_intf_10.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_10.quit_loop_state0 = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3344.ap_ST_fsm_state2;
    assign seq_loop_intf_10.quit_states_valid = 1'b1;
    assign seq_loop_intf_10.cur_state = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3344.ap_CS_fsm;
    assign seq_loop_intf_10.iter_start_state = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3344.ap_ST_fsm_state2;
    assign seq_loop_intf_10.iter_end_state0 = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3344.ap_ST_fsm_state4;
    assign seq_loop_intf_10.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_10.one_state_loop = 1'b0;
    assign seq_loop_intf_10.one_state_block = 1'b0;
    assign seq_loop_intf_10.finish = finish;
    csv_file_dump seq_loop_csv_dumper_10;
    seq_loop_monitor #(7) seq_loop_monitor_10;
    seq_loop_intf#(7) seq_loop_intf_11(clock,reset);
    assign seq_loop_intf_11.pre_loop_state0 = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3353.ap_ST_fsm_state1;
    assign seq_loop_intf_11.pre_states_valid = 1'b1;
    assign seq_loop_intf_11.post_loop_state0 = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3353.ap_ST_fsm_state5;
    assign seq_loop_intf_11.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_11.post_loop_state1 = 7'h0;
    assign seq_loop_intf_11.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_11.quit_loop_state0 = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3353.ap_ST_fsm_state2;
    assign seq_loop_intf_11.quit_states_valid = 1'b1;
    assign seq_loop_intf_11.cur_state = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3353.ap_CS_fsm;
    assign seq_loop_intf_11.iter_start_state = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3353.ap_ST_fsm_state2;
    assign seq_loop_intf_11.iter_end_state0 = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3353.ap_ST_fsm_state4;
    assign seq_loop_intf_11.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_11.one_state_loop = 1'b0;
    assign seq_loop_intf_11.one_state_block = 1'b0;
    assign seq_loop_intf_11.finish = finish;
    csv_file_dump seq_loop_csv_dumper_11;
    seq_loop_monitor #(7) seq_loop_monitor_11;
    seq_loop_intf#(7) seq_loop_intf_12(clock,reset);
    assign seq_loop_intf_12.pre_loop_state0 = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3362.ap_ST_fsm_state1;
    assign seq_loop_intf_12.pre_states_valid = 1'b1;
    assign seq_loop_intf_12.post_loop_state0 = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3362.ap_ST_fsm_state5;
    assign seq_loop_intf_12.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_12.post_loop_state1 = 7'h0;
    assign seq_loop_intf_12.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_12.quit_loop_state0 = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3362.ap_ST_fsm_state2;
    assign seq_loop_intf_12.quit_states_valid = 1'b1;
    assign seq_loop_intf_12.cur_state = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3362.ap_CS_fsm;
    assign seq_loop_intf_12.iter_start_state = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3362.ap_ST_fsm_state2;
    assign seq_loop_intf_12.iter_end_state0 = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3362.ap_ST_fsm_state4;
    assign seq_loop_intf_12.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_12.one_state_loop = 1'b0;
    assign seq_loop_intf_12.one_state_block = 1'b0;
    assign seq_loop_intf_12.finish = finish;
    csv_file_dump seq_loop_csv_dumper_12;
    seq_loop_monitor #(7) seq_loop_monitor_12;
    seq_loop_intf#(16) seq_loop_intf_13(clock,reset);
    assign seq_loop_intf_13.pre_loop_state0 = AESL_inst_TOP.grp_KBEST_fu_461.ap_ST_fsm_state5;
    assign seq_loop_intf_13.pre_states_valid = 1'b1;
    assign seq_loop_intf_13.post_loop_state0 = AESL_inst_TOP.grp_KBEST_fu_461.ap_ST_fsm_state12;
    assign seq_loop_intf_13.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_13.post_loop_state1 = AESL_inst_TOP.grp_KBEST_fu_461.ap_ST_fsm_state13;
    assign seq_loop_intf_13.post_states_valid[1] = 1'b1;
    assign seq_loop_intf_13.quit_loop_state0 = AESL_inst_TOP.grp_KBEST_fu_461.ap_ST_fsm_state6;
    assign seq_loop_intf_13.quit_states_valid = 1'b1;
    assign seq_loop_intf_13.cur_state = AESL_inst_TOP.grp_KBEST_fu_461.ap_CS_fsm;
    assign seq_loop_intf_13.iter_start_state = AESL_inst_TOP.grp_KBEST_fu_461.ap_ST_fsm_state6;
    assign seq_loop_intf_13.iter_end_state0 = AESL_inst_TOP.grp_KBEST_fu_461.ap_ST_fsm_state11;
    assign seq_loop_intf_13.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_13.one_state_loop = 1'b0;
    assign seq_loop_intf_13.one_state_block = 1'b0;
    assign seq_loop_intf_13.finish = finish;
    csv_file_dump seq_loop_csv_dumper_13;
    seq_loop_monitor #(16) seq_loop_monitor_13;
    seq_loop_intf#(16) seq_loop_intf_14(clock,reset);
    assign seq_loop_intf_14.pre_loop_state0 = AESL_inst_TOP.grp_KBEST_fu_461.ap_ST_fsm_state2;
    assign seq_loop_intf_14.pre_states_valid = 1'b1;
    assign seq_loop_intf_14.post_loop_state0 = AESL_inst_TOP.grp_KBEST_fu_461.ap_ST_fsm_state16;
    assign seq_loop_intf_14.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_14.post_loop_state1 = 16'h0;
    assign seq_loop_intf_14.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_14.quit_loop_state0 = AESL_inst_TOP.grp_KBEST_fu_461.ap_ST_fsm_state3;
    assign seq_loop_intf_14.quit_states_valid = 1'b1;
    assign seq_loop_intf_14.cur_state = AESL_inst_TOP.grp_KBEST_fu_461.ap_CS_fsm;
    assign seq_loop_intf_14.iter_start_state = AESL_inst_TOP.grp_KBEST_fu_461.ap_ST_fsm_state3;
    assign seq_loop_intf_14.iter_end_state0 = AESL_inst_TOP.grp_KBEST_fu_461.ap_ST_fsm_state15;
    assign seq_loop_intf_14.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_14.one_state_loop = 1'b0;
    assign seq_loop_intf_14.one_state_block = 1'b0;
    assign seq_loop_intf_14.finish = finish;
    csv_file_dump seq_loop_csv_dumper_14;
    seq_loop_monitor #(16) seq_loop_monitor_14;
    upc_loop_intf#(1) upc_loop_intf_1(clock,reset);
    assign upc_loop_intf_1.cur_state = AESL_inst_TOP.grp_Rayleigh_fu_311.grp_seedInitialization_fu_40.grp_seedInitialization_Pipeline_SEED_INIT_LOOP_fu_94.ap_CS_fsm;
    assign upc_loop_intf_1.iter_start_state = AESL_inst_TOP.grp_Rayleigh_fu_311.grp_seedInitialization_fu_40.grp_seedInitialization_Pipeline_SEED_INIT_LOOP_fu_94.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_1.iter_end_state = AESL_inst_TOP.grp_Rayleigh_fu_311.grp_seedInitialization_fu_40.grp_seedInitialization_Pipeline_SEED_INIT_LOOP_fu_94.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_1.quit_state = AESL_inst_TOP.grp_Rayleigh_fu_311.grp_seedInitialization_fu_40.grp_seedInitialization_Pipeline_SEED_INIT_LOOP_fu_94.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_1.iter_start_block = AESL_inst_TOP.grp_Rayleigh_fu_311.grp_seedInitialization_fu_40.grp_seedInitialization_Pipeline_SEED_INIT_LOOP_fu_94.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_1.iter_end_block = AESL_inst_TOP.grp_Rayleigh_fu_311.grp_seedInitialization_fu_40.grp_seedInitialization_Pipeline_SEED_INIT_LOOP_fu_94.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_1.quit_block = AESL_inst_TOP.grp_Rayleigh_fu_311.grp_seedInitialization_fu_40.grp_seedInitialization_Pipeline_SEED_INIT_LOOP_fu_94.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_1.iter_start_enable = AESL_inst_TOP.grp_Rayleigh_fu_311.grp_seedInitialization_fu_40.grp_seedInitialization_Pipeline_SEED_INIT_LOOP_fu_94.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_1.iter_end_enable = AESL_inst_TOP.grp_Rayleigh_fu_311.grp_seedInitialization_fu_40.grp_seedInitialization_Pipeline_SEED_INIT_LOOP_fu_94.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_1.quit_enable = AESL_inst_TOP.grp_Rayleigh_fu_311.grp_seedInitialization_fu_40.grp_seedInitialization_Pipeline_SEED_INIT_LOOP_fu_94.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_1.loop_start = AESL_inst_TOP.grp_Rayleigh_fu_311.grp_seedInitialization_fu_40.grp_seedInitialization_Pipeline_SEED_INIT_LOOP_fu_94.ap_start;
    assign upc_loop_intf_1.loop_ready = AESL_inst_TOP.grp_Rayleigh_fu_311.grp_seedInitialization_fu_40.grp_seedInitialization_Pipeline_SEED_INIT_LOOP_fu_94.ap_ready;
    assign upc_loop_intf_1.loop_done = AESL_inst_TOP.grp_Rayleigh_fu_311.grp_seedInitialization_fu_40.grp_seedInitialization_Pipeline_SEED_INIT_LOOP_fu_94.ap_done_int;
    assign upc_loop_intf_1.loop_continue = 1'b1;
    assign upc_loop_intf_1.quit_at_end = 1'b1;
    assign upc_loop_intf_1.finish = finish;
    csv_file_dump upc_loop_csv_dumper_1;
    upc_loop_monitor #(1) upc_loop_monitor_1;
    upc_loop_intf#(2) upc_loop_intf_2(clock,reset);
    assign upc_loop_intf_2.cur_state = AESL_inst_TOP.grp_Rayleigh_fu_311.grp_Rayleigh_Pipeline_VITIS_LOOP_28_1_VITIS_LOOP_29_2_fu_54.ap_CS_fsm;
    assign upc_loop_intf_2.iter_start_state = AESL_inst_TOP.grp_Rayleigh_fu_311.grp_Rayleigh_Pipeline_VITIS_LOOP_28_1_VITIS_LOOP_29_2_fu_54.ap_ST_fsm_pp0_stage1;
    assign upc_loop_intf_2.iter_end_state = AESL_inst_TOP.grp_Rayleigh_fu_311.grp_Rayleigh_Pipeline_VITIS_LOOP_28_1_VITIS_LOOP_29_2_fu_54.ap_ST_fsm_pp0_stage1;
    assign upc_loop_intf_2.quit_state = AESL_inst_TOP.grp_Rayleigh_fu_311.grp_Rayleigh_Pipeline_VITIS_LOOP_28_1_VITIS_LOOP_29_2_fu_54.ap_ST_fsm_pp0_stage1;
    assign upc_loop_intf_2.iter_start_block = AESL_inst_TOP.grp_Rayleigh_fu_311.grp_Rayleigh_Pipeline_VITIS_LOOP_28_1_VITIS_LOOP_29_2_fu_54.ap_block_pp0_stage1_subdone;
    assign upc_loop_intf_2.iter_end_block = AESL_inst_TOP.grp_Rayleigh_fu_311.grp_Rayleigh_Pipeline_VITIS_LOOP_28_1_VITIS_LOOP_29_2_fu_54.ap_block_pp0_stage1_subdone;
    assign upc_loop_intf_2.quit_block = AESL_inst_TOP.grp_Rayleigh_fu_311.grp_Rayleigh_Pipeline_VITIS_LOOP_28_1_VITIS_LOOP_29_2_fu_54.ap_block_pp0_stage1_subdone;
    assign upc_loop_intf_2.iter_start_enable = AESL_inst_TOP.grp_Rayleigh_fu_311.grp_Rayleigh_Pipeline_VITIS_LOOP_28_1_VITIS_LOOP_29_2_fu_54.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_2.iter_end_enable = AESL_inst_TOP.grp_Rayleigh_fu_311.grp_Rayleigh_Pipeline_VITIS_LOOP_28_1_VITIS_LOOP_29_2_fu_54.ap_enable_reg_pp0_iter14;
    assign upc_loop_intf_2.quit_enable = AESL_inst_TOP.grp_Rayleigh_fu_311.grp_Rayleigh_Pipeline_VITIS_LOOP_28_1_VITIS_LOOP_29_2_fu_54.ap_enable_reg_pp0_iter14;
    assign upc_loop_intf_2.loop_start = AESL_inst_TOP.grp_Rayleigh_fu_311.grp_Rayleigh_Pipeline_VITIS_LOOP_28_1_VITIS_LOOP_29_2_fu_54.ap_start;
    assign upc_loop_intf_2.loop_ready = AESL_inst_TOP.grp_Rayleigh_fu_311.grp_Rayleigh_Pipeline_VITIS_LOOP_28_1_VITIS_LOOP_29_2_fu_54.ap_ready;
    assign upc_loop_intf_2.loop_done = AESL_inst_TOP.grp_Rayleigh_fu_311.grp_Rayleigh_Pipeline_VITIS_LOOP_28_1_VITIS_LOOP_29_2_fu_54.ap_done_int;
    assign upc_loop_intf_2.loop_continue = 1'b1;
    assign upc_loop_intf_2.quit_at_end = 1'b1;
    assign upc_loop_intf_2.finish = finish;
    csv_file_dump upc_loop_csv_dumper_2;
    upc_loop_monitor #(2) upc_loop_monitor_2;
    upc_loop_intf#(2) upc_loop_intf_3(clock,reset);
    assign upc_loop_intf_3.cur_state = AESL_inst_TOP.grp_Rayleigh_fu_311.grp_Rayleigh_Pipeline_VITIS_LOOP_40_3_VITIS_LOOP_41_4_fu_66.ap_CS_fsm;
    assign upc_loop_intf_3.iter_start_state = AESL_inst_TOP.grp_Rayleigh_fu_311.grp_Rayleigh_Pipeline_VITIS_LOOP_40_3_VITIS_LOOP_41_4_fu_66.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_3.iter_end_state = AESL_inst_TOP.grp_Rayleigh_fu_311.grp_Rayleigh_Pipeline_VITIS_LOOP_40_3_VITIS_LOOP_41_4_fu_66.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_3.quit_state = AESL_inst_TOP.grp_Rayleigh_fu_311.grp_Rayleigh_Pipeline_VITIS_LOOP_40_3_VITIS_LOOP_41_4_fu_66.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_3.iter_start_block = AESL_inst_TOP.grp_Rayleigh_fu_311.grp_Rayleigh_Pipeline_VITIS_LOOP_40_3_VITIS_LOOP_41_4_fu_66.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_3.iter_end_block = AESL_inst_TOP.grp_Rayleigh_fu_311.grp_Rayleigh_Pipeline_VITIS_LOOP_40_3_VITIS_LOOP_41_4_fu_66.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_3.quit_block = AESL_inst_TOP.grp_Rayleigh_fu_311.grp_Rayleigh_Pipeline_VITIS_LOOP_40_3_VITIS_LOOP_41_4_fu_66.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_3.iter_start_enable = AESL_inst_TOP.grp_Rayleigh_fu_311.grp_Rayleigh_Pipeline_VITIS_LOOP_40_3_VITIS_LOOP_41_4_fu_66.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_3.iter_end_enable = AESL_inst_TOP.grp_Rayleigh_fu_311.grp_Rayleigh_Pipeline_VITIS_LOOP_40_3_VITIS_LOOP_41_4_fu_66.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_3.quit_enable = AESL_inst_TOP.grp_Rayleigh_fu_311.grp_Rayleigh_Pipeline_VITIS_LOOP_40_3_VITIS_LOOP_41_4_fu_66.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_3.loop_start = AESL_inst_TOP.grp_Rayleigh_fu_311.grp_Rayleigh_Pipeline_VITIS_LOOP_40_3_VITIS_LOOP_41_4_fu_66.ap_start;
    assign upc_loop_intf_3.loop_ready = AESL_inst_TOP.grp_Rayleigh_fu_311.grp_Rayleigh_Pipeline_VITIS_LOOP_40_3_VITIS_LOOP_41_4_fu_66.ap_ready;
    assign upc_loop_intf_3.loop_done = AESL_inst_TOP.grp_Rayleigh_fu_311.grp_Rayleigh_Pipeline_VITIS_LOOP_40_3_VITIS_LOOP_41_4_fu_66.ap_done_int;
    assign upc_loop_intf_3.loop_continue = 1'b1;
    assign upc_loop_intf_3.quit_at_end = 1'b0;
    assign upc_loop_intf_3.finish = finish;
    csv_file_dump upc_loop_csv_dumper_3;
    upc_loop_monitor #(2) upc_loop_monitor_3;
    upc_loop_intf#(4) upc_loop_intf_4(clock,reset);
    assign upc_loop_intf_4.cur_state = AESL_inst_TOP.grp_Rayleigh_fu_311.grp_Rayleigh_Pipeline_VITIS_LOOP_69_6_fu_74.ap_CS_fsm;
    assign upc_loop_intf_4.iter_start_state = AESL_inst_TOP.grp_Rayleigh_fu_311.grp_Rayleigh_Pipeline_VITIS_LOOP_69_6_fu_74.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_4.iter_end_state = AESL_inst_TOP.grp_Rayleigh_fu_311.grp_Rayleigh_Pipeline_VITIS_LOOP_69_6_fu_74.ap_ST_fsm_pp0_stage1;
    assign upc_loop_intf_4.quit_state = AESL_inst_TOP.grp_Rayleigh_fu_311.grp_Rayleigh_Pipeline_VITIS_LOOP_69_6_fu_74.ap_ST_fsm_pp0_stage1;
    assign upc_loop_intf_4.iter_start_block = AESL_inst_TOP.grp_Rayleigh_fu_311.grp_Rayleigh_Pipeline_VITIS_LOOP_69_6_fu_74.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_4.iter_end_block = AESL_inst_TOP.grp_Rayleigh_fu_311.grp_Rayleigh_Pipeline_VITIS_LOOP_69_6_fu_74.ap_block_pp0_stage1_subdone;
    assign upc_loop_intf_4.quit_block = AESL_inst_TOP.grp_Rayleigh_fu_311.grp_Rayleigh_Pipeline_VITIS_LOOP_69_6_fu_74.ap_block_pp0_stage1_subdone;
    assign upc_loop_intf_4.iter_start_enable = AESL_inst_TOP.grp_Rayleigh_fu_311.grp_Rayleigh_Pipeline_VITIS_LOOP_69_6_fu_74.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_4.iter_end_enable = AESL_inst_TOP.grp_Rayleigh_fu_311.grp_Rayleigh_Pipeline_VITIS_LOOP_69_6_fu_74.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_4.quit_enable = AESL_inst_TOP.grp_Rayleigh_fu_311.grp_Rayleigh_Pipeline_VITIS_LOOP_69_6_fu_74.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_4.loop_start = AESL_inst_TOP.grp_Rayleigh_fu_311.grp_Rayleigh_Pipeline_VITIS_LOOP_69_6_fu_74.ap_start;
    assign upc_loop_intf_4.loop_ready = AESL_inst_TOP.grp_Rayleigh_fu_311.grp_Rayleigh_Pipeline_VITIS_LOOP_69_6_fu_74.ap_ready;
    assign upc_loop_intf_4.loop_done = AESL_inst_TOP.grp_Rayleigh_fu_311.grp_Rayleigh_Pipeline_VITIS_LOOP_69_6_fu_74.ap_done_int;
    assign upc_loop_intf_4.loop_continue = 1'b1;
    assign upc_loop_intf_4.quit_at_end = 1'b1;
    assign upc_loop_intf_4.finish = finish;
    csv_file_dump upc_loop_csv_dumper_4;
    upc_loop_monitor #(4) upc_loop_monitor_4;
    upc_loop_intf#(1) upc_loop_intf_5(clock,reset);
    assign upc_loop_intf_5.cur_state = AESL_inst_TOP.grp_AWGN_fu_319.grp_seedInitialization_fu_432.grp_seedInitialization_Pipeline_SEED_INIT_LOOP_fu_94.ap_CS_fsm;
    assign upc_loop_intf_5.iter_start_state = AESL_inst_TOP.grp_AWGN_fu_319.grp_seedInitialization_fu_432.grp_seedInitialization_Pipeline_SEED_INIT_LOOP_fu_94.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_5.iter_end_state = AESL_inst_TOP.grp_AWGN_fu_319.grp_seedInitialization_fu_432.grp_seedInitialization_Pipeline_SEED_INIT_LOOP_fu_94.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_5.quit_state = AESL_inst_TOP.grp_AWGN_fu_319.grp_seedInitialization_fu_432.grp_seedInitialization_Pipeline_SEED_INIT_LOOP_fu_94.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_5.iter_start_block = AESL_inst_TOP.grp_AWGN_fu_319.grp_seedInitialization_fu_432.grp_seedInitialization_Pipeline_SEED_INIT_LOOP_fu_94.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_5.iter_end_block = AESL_inst_TOP.grp_AWGN_fu_319.grp_seedInitialization_fu_432.grp_seedInitialization_Pipeline_SEED_INIT_LOOP_fu_94.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_5.quit_block = AESL_inst_TOP.grp_AWGN_fu_319.grp_seedInitialization_fu_432.grp_seedInitialization_Pipeline_SEED_INIT_LOOP_fu_94.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_5.iter_start_enable = AESL_inst_TOP.grp_AWGN_fu_319.grp_seedInitialization_fu_432.grp_seedInitialization_Pipeline_SEED_INIT_LOOP_fu_94.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_5.iter_end_enable = AESL_inst_TOP.grp_AWGN_fu_319.grp_seedInitialization_fu_432.grp_seedInitialization_Pipeline_SEED_INIT_LOOP_fu_94.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_5.quit_enable = AESL_inst_TOP.grp_AWGN_fu_319.grp_seedInitialization_fu_432.grp_seedInitialization_Pipeline_SEED_INIT_LOOP_fu_94.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_5.loop_start = AESL_inst_TOP.grp_AWGN_fu_319.grp_seedInitialization_fu_432.grp_seedInitialization_Pipeline_SEED_INIT_LOOP_fu_94.ap_start;
    assign upc_loop_intf_5.loop_ready = AESL_inst_TOP.grp_AWGN_fu_319.grp_seedInitialization_fu_432.grp_seedInitialization_Pipeline_SEED_INIT_LOOP_fu_94.ap_ready;
    assign upc_loop_intf_5.loop_done = AESL_inst_TOP.grp_AWGN_fu_319.grp_seedInitialization_fu_432.grp_seedInitialization_Pipeline_SEED_INIT_LOOP_fu_94.ap_done_int;
    assign upc_loop_intf_5.loop_continue = 1'b1;
    assign upc_loop_intf_5.quit_at_end = 1'b1;
    assign upc_loop_intf_5.finish = finish;
    csv_file_dump upc_loop_csv_dumper_5;
    upc_loop_monitor #(1) upc_loop_monitor_5;
    upc_loop_intf#(1) upc_loop_intf_6(clock,reset);
    assign upc_loop_intf_6.cur_state = AESL_inst_TOP.grp_TOP_Pipeline_VITIS_LOOP_482_2_VITIS_LOOP_483_3_fu_325.ap_CS_fsm;
    assign upc_loop_intf_6.iter_start_state = AESL_inst_TOP.grp_TOP_Pipeline_VITIS_LOOP_482_2_VITIS_LOOP_483_3_fu_325.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_6.iter_end_state = AESL_inst_TOP.grp_TOP_Pipeline_VITIS_LOOP_482_2_VITIS_LOOP_483_3_fu_325.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_6.quit_state = AESL_inst_TOP.grp_TOP_Pipeline_VITIS_LOOP_482_2_VITIS_LOOP_483_3_fu_325.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_6.iter_start_block = AESL_inst_TOP.grp_TOP_Pipeline_VITIS_LOOP_482_2_VITIS_LOOP_483_3_fu_325.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_6.iter_end_block = AESL_inst_TOP.grp_TOP_Pipeline_VITIS_LOOP_482_2_VITIS_LOOP_483_3_fu_325.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_6.quit_block = AESL_inst_TOP.grp_TOP_Pipeline_VITIS_LOOP_482_2_VITIS_LOOP_483_3_fu_325.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_6.iter_start_enable = AESL_inst_TOP.grp_TOP_Pipeline_VITIS_LOOP_482_2_VITIS_LOOP_483_3_fu_325.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_6.iter_end_enable = AESL_inst_TOP.grp_TOP_Pipeline_VITIS_LOOP_482_2_VITIS_LOOP_483_3_fu_325.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_6.quit_enable = AESL_inst_TOP.grp_TOP_Pipeline_VITIS_LOOP_482_2_VITIS_LOOP_483_3_fu_325.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_6.loop_start = AESL_inst_TOP.grp_TOP_Pipeline_VITIS_LOOP_482_2_VITIS_LOOP_483_3_fu_325.ap_start;
    assign upc_loop_intf_6.loop_ready = AESL_inst_TOP.grp_TOP_Pipeline_VITIS_LOOP_482_2_VITIS_LOOP_483_3_fu_325.ap_ready;
    assign upc_loop_intf_6.loop_done = AESL_inst_TOP.grp_TOP_Pipeline_VITIS_LOOP_482_2_VITIS_LOOP_483_3_fu_325.ap_done_int;
    assign upc_loop_intf_6.loop_continue = 1'b1;
    assign upc_loop_intf_6.quit_at_end = 1'b0;
    assign upc_loop_intf_6.finish = finish;
    csv_file_dump upc_loop_csv_dumper_6;
    upc_loop_monitor #(1) upc_loop_monitor_6;
    upc_loop_intf#(1) upc_loop_intf_7(clock,reset);
    assign upc_loop_intf_7.cur_state = AESL_inst_TOP.grp_TOP_Pipeline_VITIS_LOOP_488_4_fu_346.ap_CS_fsm;
    assign upc_loop_intf_7.iter_start_state = AESL_inst_TOP.grp_TOP_Pipeline_VITIS_LOOP_488_4_fu_346.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_7.iter_end_state = AESL_inst_TOP.grp_TOP_Pipeline_VITIS_LOOP_488_4_fu_346.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_7.quit_state = AESL_inst_TOP.grp_TOP_Pipeline_VITIS_LOOP_488_4_fu_346.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_7.iter_start_block = AESL_inst_TOP.grp_TOP_Pipeline_VITIS_LOOP_488_4_fu_346.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_7.iter_end_block = AESL_inst_TOP.grp_TOP_Pipeline_VITIS_LOOP_488_4_fu_346.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_7.quit_block = AESL_inst_TOP.grp_TOP_Pipeline_VITIS_LOOP_488_4_fu_346.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_7.iter_start_enable = AESL_inst_TOP.grp_TOP_Pipeline_VITIS_LOOP_488_4_fu_346.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_7.iter_end_enable = AESL_inst_TOP.grp_TOP_Pipeline_VITIS_LOOP_488_4_fu_346.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_7.quit_enable = AESL_inst_TOP.grp_TOP_Pipeline_VITIS_LOOP_488_4_fu_346.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_7.loop_start = AESL_inst_TOP.grp_TOP_Pipeline_VITIS_LOOP_488_4_fu_346.ap_start;
    assign upc_loop_intf_7.loop_ready = AESL_inst_TOP.grp_TOP_Pipeline_VITIS_LOOP_488_4_fu_346.ap_ready;
    assign upc_loop_intf_7.loop_done = AESL_inst_TOP.grp_TOP_Pipeline_VITIS_LOOP_488_4_fu_346.ap_done_int;
    assign upc_loop_intf_7.loop_continue = 1'b1;
    assign upc_loop_intf_7.quit_at_end = 1'b0;
    assign upc_loop_intf_7.finish = finish;
    csv_file_dump upc_loop_csv_dumper_7;
    upc_loop_monitor #(1) upc_loop_monitor_7;
    upc_loop_intf#(1) upc_loop_intf_8(clock,reset);
    assign upc_loop_intf_8.cur_state = AESL_inst_TOP.grp_TOP_Pipeline_VITIS_LOOP_492_5_VITIS_LOOP_493_6_fu_352.ap_CS_fsm;
    assign upc_loop_intf_8.iter_start_state = AESL_inst_TOP.grp_TOP_Pipeline_VITIS_LOOP_492_5_VITIS_LOOP_493_6_fu_352.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_8.iter_end_state = AESL_inst_TOP.grp_TOP_Pipeline_VITIS_LOOP_492_5_VITIS_LOOP_493_6_fu_352.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_8.quit_state = AESL_inst_TOP.grp_TOP_Pipeline_VITIS_LOOP_492_5_VITIS_LOOP_493_6_fu_352.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_8.iter_start_block = AESL_inst_TOP.grp_TOP_Pipeline_VITIS_LOOP_492_5_VITIS_LOOP_493_6_fu_352.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_8.iter_end_block = AESL_inst_TOP.grp_TOP_Pipeline_VITIS_LOOP_492_5_VITIS_LOOP_493_6_fu_352.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_8.quit_block = AESL_inst_TOP.grp_TOP_Pipeline_VITIS_LOOP_492_5_VITIS_LOOP_493_6_fu_352.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_8.iter_start_enable = AESL_inst_TOP.grp_TOP_Pipeline_VITIS_LOOP_492_5_VITIS_LOOP_493_6_fu_352.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_8.iter_end_enable = AESL_inst_TOP.grp_TOP_Pipeline_VITIS_LOOP_492_5_VITIS_LOOP_493_6_fu_352.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_8.quit_enable = AESL_inst_TOP.grp_TOP_Pipeline_VITIS_LOOP_492_5_VITIS_LOOP_493_6_fu_352.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_8.loop_start = AESL_inst_TOP.grp_TOP_Pipeline_VITIS_LOOP_492_5_VITIS_LOOP_493_6_fu_352.ap_start;
    assign upc_loop_intf_8.loop_ready = AESL_inst_TOP.grp_TOP_Pipeline_VITIS_LOOP_492_5_VITIS_LOOP_493_6_fu_352.ap_ready;
    assign upc_loop_intf_8.loop_done = AESL_inst_TOP.grp_TOP_Pipeline_VITIS_LOOP_492_5_VITIS_LOOP_493_6_fu_352.ap_done_int;
    assign upc_loop_intf_8.loop_continue = 1'b1;
    assign upc_loop_intf_8.quit_at_end = 1'b0;
    assign upc_loop_intf_8.finish = finish;
    csv_file_dump upc_loop_csv_dumper_8;
    upc_loop_monitor #(1) upc_loop_monitor_8;
    upc_loop_intf#(1) upc_loop_intf_9(clock,reset);
    assign upc_loop_intf_9.cur_state = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_V_fu_3293.grp_CORDIC_V_Pipeline_VITIS_LOOP_94_2_fu_173.ap_CS_fsm;
    assign upc_loop_intf_9.iter_start_state = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_V_fu_3293.grp_CORDIC_V_Pipeline_VITIS_LOOP_94_2_fu_173.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_9.iter_end_state = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_V_fu_3293.grp_CORDIC_V_Pipeline_VITIS_LOOP_94_2_fu_173.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_9.quit_state = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_V_fu_3293.grp_CORDIC_V_Pipeline_VITIS_LOOP_94_2_fu_173.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_9.iter_start_block = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_V_fu_3293.grp_CORDIC_V_Pipeline_VITIS_LOOP_94_2_fu_173.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_9.iter_end_block = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_V_fu_3293.grp_CORDIC_V_Pipeline_VITIS_LOOP_94_2_fu_173.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_9.quit_block = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_V_fu_3293.grp_CORDIC_V_Pipeline_VITIS_LOOP_94_2_fu_173.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_9.iter_start_enable = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_V_fu_3293.grp_CORDIC_V_Pipeline_VITIS_LOOP_94_2_fu_173.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_9.iter_end_enable = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_V_fu_3293.grp_CORDIC_V_Pipeline_VITIS_LOOP_94_2_fu_173.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_9.quit_enable = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_V_fu_3293.grp_CORDIC_V_Pipeline_VITIS_LOOP_94_2_fu_173.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_9.loop_start = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_V_fu_3293.grp_CORDIC_V_Pipeline_VITIS_LOOP_94_2_fu_173.ap_start;
    assign upc_loop_intf_9.loop_ready = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_V_fu_3293.grp_CORDIC_V_Pipeline_VITIS_LOOP_94_2_fu_173.ap_ready;
    assign upc_loop_intf_9.loop_done = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_V_fu_3293.grp_CORDIC_V_Pipeline_VITIS_LOOP_94_2_fu_173.ap_done_int;
    assign upc_loop_intf_9.loop_continue = 1'b1;
    assign upc_loop_intf_9.quit_at_end = 1'b1;
    assign upc_loop_intf_9.finish = finish;
    csv_file_dump upc_loop_csv_dumper_9;
    upc_loop_monitor #(1) upc_loop_monitor_9;
    upc_loop_intf#(1) upc_loop_intf_10(clock,reset);
    assign upc_loop_intf_10.cur_state = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3308.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_CS_fsm;
    assign upc_loop_intf_10.iter_start_state = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3308.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_10.iter_end_state = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3308.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_10.quit_state = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3308.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_10.iter_start_block = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3308.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_10.iter_end_block = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3308.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_10.quit_block = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3308.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_10.iter_start_enable = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3308.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_10.iter_end_enable = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3308.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_10.quit_enable = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3308.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_10.loop_start = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3308.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_start;
    assign upc_loop_intf_10.loop_ready = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3308.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_ready;
    assign upc_loop_intf_10.loop_done = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3308.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_done_int;
    assign upc_loop_intf_10.loop_continue = 1'b1;
    assign upc_loop_intf_10.quit_at_end = 1'b1;
    assign upc_loop_intf_10.finish = finish;
    csv_file_dump upc_loop_csv_dumper_10;
    upc_loop_monitor #(1) upc_loop_monitor_10;
    upc_loop_intf#(1) upc_loop_intf_11(clock,reset);
    assign upc_loop_intf_11.cur_state = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3326.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_CS_fsm;
    assign upc_loop_intf_11.iter_start_state = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3326.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_11.iter_end_state = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3326.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_11.quit_state = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3326.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_11.iter_start_block = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3326.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_11.iter_end_block = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3326.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_11.quit_block = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3326.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_11.iter_start_enable = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3326.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_11.iter_end_enable = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3326.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_11.quit_enable = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3326.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_11.loop_start = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3326.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_start;
    assign upc_loop_intf_11.loop_ready = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3326.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_ready;
    assign upc_loop_intf_11.loop_done = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3326.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_done_int;
    assign upc_loop_intf_11.loop_continue = 1'b1;
    assign upc_loop_intf_11.quit_at_end = 1'b1;
    assign upc_loop_intf_11.finish = finish;
    csv_file_dump upc_loop_csv_dumper_11;
    upc_loop_monitor #(1) upc_loop_monitor_11;
    upc_loop_intf#(1) upc_loop_intf_12(clock,reset);
    assign upc_loop_intf_12.cur_state = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3335.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_CS_fsm;
    assign upc_loop_intf_12.iter_start_state = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3335.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_12.iter_end_state = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3335.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_12.quit_state = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3335.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_12.iter_start_block = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3335.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_12.iter_end_block = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3335.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_12.quit_block = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3335.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_12.iter_start_enable = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3335.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_12.iter_end_enable = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3335.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_12.quit_enable = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3335.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_12.loop_start = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3335.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_start;
    assign upc_loop_intf_12.loop_ready = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3335.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_ready;
    assign upc_loop_intf_12.loop_done = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3335.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_done_int;
    assign upc_loop_intf_12.loop_continue = 1'b1;
    assign upc_loop_intf_12.quit_at_end = 1'b1;
    assign upc_loop_intf_12.finish = finish;
    csv_file_dump upc_loop_csv_dumper_12;
    upc_loop_monitor #(1) upc_loop_monitor_12;
    upc_loop_intf#(1) upc_loop_intf_13(clock,reset);
    assign upc_loop_intf_13.cur_state = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3344.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_CS_fsm;
    assign upc_loop_intf_13.iter_start_state = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3344.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_13.iter_end_state = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3344.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_13.quit_state = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3344.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_13.iter_start_block = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3344.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_13.iter_end_block = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3344.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_13.quit_block = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3344.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_13.iter_start_enable = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3344.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_13.iter_end_enable = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3344.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_13.quit_enable = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3344.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_13.loop_start = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3344.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_start;
    assign upc_loop_intf_13.loop_ready = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3344.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_ready;
    assign upc_loop_intf_13.loop_done = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3344.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_done_int;
    assign upc_loop_intf_13.loop_continue = 1'b1;
    assign upc_loop_intf_13.quit_at_end = 1'b1;
    assign upc_loop_intf_13.finish = finish;
    csv_file_dump upc_loop_csv_dumper_13;
    upc_loop_monitor #(1) upc_loop_monitor_13;
    upc_loop_intf#(1) upc_loop_intf_14(clock,reset);
    assign upc_loop_intf_14.cur_state = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3353.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_CS_fsm;
    assign upc_loop_intf_14.iter_start_state = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3353.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_14.iter_end_state = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3353.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_14.quit_state = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3353.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_14.iter_start_block = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3353.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_14.iter_end_block = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3353.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_14.quit_block = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3353.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_14.iter_start_enable = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3353.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_14.iter_end_enable = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3353.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_14.quit_enable = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3353.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_14.loop_start = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3353.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_start;
    assign upc_loop_intf_14.loop_ready = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3353.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_ready;
    assign upc_loop_intf_14.loop_done = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3353.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_done_int;
    assign upc_loop_intf_14.loop_continue = 1'b1;
    assign upc_loop_intf_14.quit_at_end = 1'b1;
    assign upc_loop_intf_14.finish = finish;
    csv_file_dump upc_loop_csv_dumper_14;
    upc_loop_monitor #(1) upc_loop_monitor_14;
    upc_loop_intf#(1) upc_loop_intf_15(clock,reset);
    assign upc_loop_intf_15.cur_state = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3362.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_CS_fsm;
    assign upc_loop_intf_15.iter_start_state = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3362.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_15.iter_end_state = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3362.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_15.quit_state = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3362.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_15.iter_start_block = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3362.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_15.iter_end_block = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3362.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_15.quit_block = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3362.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_15.iter_start_enable = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3362.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_15.iter_end_enable = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3362.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_15.quit_enable = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3362.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_15.loop_start = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3362.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_start;
    assign upc_loop_intf_15.loop_ready = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3362.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_ready;
    assign upc_loop_intf_15.loop_done = AESL_inst_TOP.grp_QRD_fu_389.grp_CORDIC_R_fu_3362.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_157.ap_done_int;
    assign upc_loop_intf_15.loop_continue = 1'b1;
    assign upc_loop_intf_15.quit_at_end = 1'b1;
    assign upc_loop_intf_15.finish = finish;
    csv_file_dump upc_loop_csv_dumper_15;
    upc_loop_monitor #(1) upc_loop_monitor_15;
    upc_loop_intf#(27) upc_loop_intf_16(clock,reset);
    assign upc_loop_intf_16.cur_state = AESL_inst_TOP.grp_QRD_fu_389.grp_QRD_Pipeline_VITIS_LOOP_268_8_fu_3539.ap_CS_fsm;
    assign upc_loop_intf_16.iter_start_state = AESL_inst_TOP.grp_QRD_fu_389.grp_QRD_Pipeline_VITIS_LOOP_268_8_fu_3539.ap_ST_fsm_pp0_stage1;
    assign upc_loop_intf_16.iter_end_state = AESL_inst_TOP.grp_QRD_fu_389.grp_QRD_Pipeline_VITIS_LOOP_268_8_fu_3539.ap_ST_fsm_pp0_stage1;
    assign upc_loop_intf_16.quit_state = AESL_inst_TOP.grp_QRD_fu_389.grp_QRD_Pipeline_VITIS_LOOP_268_8_fu_3539.ap_ST_fsm_pp0_stage1;
    assign upc_loop_intf_16.iter_start_block = AESL_inst_TOP.grp_QRD_fu_389.grp_QRD_Pipeline_VITIS_LOOP_268_8_fu_3539.ap_block_pp0_stage1_subdone;
    assign upc_loop_intf_16.iter_end_block = AESL_inst_TOP.grp_QRD_fu_389.grp_QRD_Pipeline_VITIS_LOOP_268_8_fu_3539.ap_block_pp0_stage1_subdone;
    assign upc_loop_intf_16.quit_block = AESL_inst_TOP.grp_QRD_fu_389.grp_QRD_Pipeline_VITIS_LOOP_268_8_fu_3539.ap_block_pp0_stage1_subdone;
    assign upc_loop_intf_16.iter_start_enable = AESL_inst_TOP.grp_QRD_fu_389.grp_QRD_Pipeline_VITIS_LOOP_268_8_fu_3539.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_16.iter_end_enable = AESL_inst_TOP.grp_QRD_fu_389.grp_QRD_Pipeline_VITIS_LOOP_268_8_fu_3539.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_16.quit_enable = AESL_inst_TOP.grp_QRD_fu_389.grp_QRD_Pipeline_VITIS_LOOP_268_8_fu_3539.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_16.loop_start = AESL_inst_TOP.grp_QRD_fu_389.grp_QRD_Pipeline_VITIS_LOOP_268_8_fu_3539.ap_start;
    assign upc_loop_intf_16.loop_ready = AESL_inst_TOP.grp_QRD_fu_389.grp_QRD_Pipeline_VITIS_LOOP_268_8_fu_3539.ap_ready;
    assign upc_loop_intf_16.loop_done = AESL_inst_TOP.grp_QRD_fu_389.grp_QRD_Pipeline_VITIS_LOOP_268_8_fu_3539.ap_done_int;
    assign upc_loop_intf_16.loop_continue = 1'b1;
    assign upc_loop_intf_16.quit_at_end = 1'b0;
    assign upc_loop_intf_16.finish = finish;
    csv_file_dump upc_loop_csv_dumper_16;
    upc_loop_monitor #(27) upc_loop_monitor_16;
    upc_loop_intf#(1) upc_loop_intf_17(clock,reset);
    assign upc_loop_intf_17.cur_state = AESL_inst_TOP.grp_QRD_fu_389.grp_QRD_Pipeline_VITIS_LOOP_316_9_VITIS_LOOP_317_10_fu_3674.ap_CS_fsm;
    assign upc_loop_intf_17.iter_start_state = AESL_inst_TOP.grp_QRD_fu_389.grp_QRD_Pipeline_VITIS_LOOP_316_9_VITIS_LOOP_317_10_fu_3674.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_17.iter_end_state = AESL_inst_TOP.grp_QRD_fu_389.grp_QRD_Pipeline_VITIS_LOOP_316_9_VITIS_LOOP_317_10_fu_3674.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_17.quit_state = AESL_inst_TOP.grp_QRD_fu_389.grp_QRD_Pipeline_VITIS_LOOP_316_9_VITIS_LOOP_317_10_fu_3674.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_17.iter_start_block = AESL_inst_TOP.grp_QRD_fu_389.grp_QRD_Pipeline_VITIS_LOOP_316_9_VITIS_LOOP_317_10_fu_3674.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_17.iter_end_block = AESL_inst_TOP.grp_QRD_fu_389.grp_QRD_Pipeline_VITIS_LOOP_316_9_VITIS_LOOP_317_10_fu_3674.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_17.quit_block = AESL_inst_TOP.grp_QRD_fu_389.grp_QRD_Pipeline_VITIS_LOOP_316_9_VITIS_LOOP_317_10_fu_3674.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_17.iter_start_enable = AESL_inst_TOP.grp_QRD_fu_389.grp_QRD_Pipeline_VITIS_LOOP_316_9_VITIS_LOOP_317_10_fu_3674.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_17.iter_end_enable = AESL_inst_TOP.grp_QRD_fu_389.grp_QRD_Pipeline_VITIS_LOOP_316_9_VITIS_LOOP_317_10_fu_3674.ap_enable_reg_pp0_iter10;
    assign upc_loop_intf_17.quit_enable = AESL_inst_TOP.grp_QRD_fu_389.grp_QRD_Pipeline_VITIS_LOOP_316_9_VITIS_LOOP_317_10_fu_3674.ap_enable_reg_pp0_iter10;
    assign upc_loop_intf_17.loop_start = AESL_inst_TOP.grp_QRD_fu_389.grp_QRD_Pipeline_VITIS_LOOP_316_9_VITIS_LOOP_317_10_fu_3674.ap_start;
    assign upc_loop_intf_17.loop_ready = AESL_inst_TOP.grp_QRD_fu_389.grp_QRD_Pipeline_VITIS_LOOP_316_9_VITIS_LOOP_317_10_fu_3674.ap_ready;
    assign upc_loop_intf_17.loop_done = AESL_inst_TOP.grp_QRD_fu_389.grp_QRD_Pipeline_VITIS_LOOP_316_9_VITIS_LOOP_317_10_fu_3674.ap_done_int;
    assign upc_loop_intf_17.loop_continue = 1'b1;
    assign upc_loop_intf_17.quit_at_end = 1'b1;
    assign upc_loop_intf_17.finish = finish;
    csv_file_dump upc_loop_csv_dumper_17;
    upc_loop_monitor #(1) upc_loop_monitor_17;
    upc_loop_intf#(1) upc_loop_intf_18(clock,reset);
    assign upc_loop_intf_18.cur_state = AESL_inst_TOP.grp_TOP_Pipeline_VITIS_LOOP_433_1_fu_445.ap_CS_fsm;
    assign upc_loop_intf_18.iter_start_state = AESL_inst_TOP.grp_TOP_Pipeline_VITIS_LOOP_433_1_fu_445.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_18.iter_end_state = AESL_inst_TOP.grp_TOP_Pipeline_VITIS_LOOP_433_1_fu_445.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_18.quit_state = AESL_inst_TOP.grp_TOP_Pipeline_VITIS_LOOP_433_1_fu_445.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_18.iter_start_block = AESL_inst_TOP.grp_TOP_Pipeline_VITIS_LOOP_433_1_fu_445.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_18.iter_end_block = AESL_inst_TOP.grp_TOP_Pipeline_VITIS_LOOP_433_1_fu_445.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_18.quit_block = AESL_inst_TOP.grp_TOP_Pipeline_VITIS_LOOP_433_1_fu_445.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_18.iter_start_enable = AESL_inst_TOP.grp_TOP_Pipeline_VITIS_LOOP_433_1_fu_445.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_18.iter_end_enable = AESL_inst_TOP.grp_TOP_Pipeline_VITIS_LOOP_433_1_fu_445.ap_enable_reg_pp0_iter11;
    assign upc_loop_intf_18.quit_enable = AESL_inst_TOP.grp_TOP_Pipeline_VITIS_LOOP_433_1_fu_445.ap_enable_reg_pp0_iter11;
    assign upc_loop_intf_18.loop_start = AESL_inst_TOP.grp_TOP_Pipeline_VITIS_LOOP_433_1_fu_445.ap_start;
    assign upc_loop_intf_18.loop_ready = AESL_inst_TOP.grp_TOP_Pipeline_VITIS_LOOP_433_1_fu_445.ap_ready;
    assign upc_loop_intf_18.loop_done = AESL_inst_TOP.grp_TOP_Pipeline_VITIS_LOOP_433_1_fu_445.ap_done_int;
    assign upc_loop_intf_18.loop_continue = 1'b1;
    assign upc_loop_intf_18.quit_at_end = 1'b1;
    assign upc_loop_intf_18.finish = finish;
    csv_file_dump upc_loop_csv_dumper_18;
    upc_loop_monitor #(1) upc_loop_monitor_18;
    upc_loop_intf#(1) upc_loop_intf_19(clock,reset);
    assign upc_loop_intf_19.cur_state = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_VITIS_LOOP_347_1_fu_939.ap_CS_fsm;
    assign upc_loop_intf_19.iter_start_state = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_VITIS_LOOP_347_1_fu_939.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_19.iter_end_state = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_VITIS_LOOP_347_1_fu_939.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_19.quit_state = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_VITIS_LOOP_347_1_fu_939.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_19.iter_start_block = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_VITIS_LOOP_347_1_fu_939.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_19.iter_end_block = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_VITIS_LOOP_347_1_fu_939.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_19.quit_block = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_VITIS_LOOP_347_1_fu_939.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_19.iter_start_enable = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_VITIS_LOOP_347_1_fu_939.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_19.iter_end_enable = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_VITIS_LOOP_347_1_fu_939.ap_enable_reg_pp0_iter4;
    assign upc_loop_intf_19.quit_enable = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_VITIS_LOOP_347_1_fu_939.ap_enable_reg_pp0_iter4;
    assign upc_loop_intf_19.loop_start = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_VITIS_LOOP_347_1_fu_939.ap_start;
    assign upc_loop_intf_19.loop_ready = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_VITIS_LOOP_347_1_fu_939.ap_ready;
    assign upc_loop_intf_19.loop_done = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_VITIS_LOOP_347_1_fu_939.ap_done_int;
    assign upc_loop_intf_19.loop_continue = 1'b1;
    assign upc_loop_intf_19.quit_at_end = 1'b1;
    assign upc_loop_intf_19.finish = finish;
    csv_file_dump upc_loop_csv_dumper_19;
    upc_loop_monitor #(1) upc_loop_monitor_19;
    upc_loop_intf#(1) upc_loop_intf_20(clock,reset);
    assign upc_loop_intf_20.cur_state = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_VITIS_LOOP_364_3_fu_947.ap_CS_fsm;
    assign upc_loop_intf_20.iter_start_state = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_VITIS_LOOP_364_3_fu_947.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_20.iter_end_state = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_VITIS_LOOP_364_3_fu_947.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_20.quit_state = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_VITIS_LOOP_364_3_fu_947.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_20.iter_start_block = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_VITIS_LOOP_364_3_fu_947.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_20.iter_end_block = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_VITIS_LOOP_364_3_fu_947.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_20.quit_block = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_VITIS_LOOP_364_3_fu_947.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_20.iter_start_enable = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_VITIS_LOOP_364_3_fu_947.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_20.iter_end_enable = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_VITIS_LOOP_364_3_fu_947.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_20.quit_enable = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_VITIS_LOOP_364_3_fu_947.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_20.loop_start = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_VITIS_LOOP_364_3_fu_947.ap_start;
    assign upc_loop_intf_20.loop_ready = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_VITIS_LOOP_364_3_fu_947.ap_ready;
    assign upc_loop_intf_20.loop_done = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_VITIS_LOOP_364_3_fu_947.ap_done_int;
    assign upc_loop_intf_20.loop_continue = 1'b1;
    assign upc_loop_intf_20.quit_at_end = 1'b0;
    assign upc_loop_intf_20.finish = finish;
    csv_file_dump upc_loop_csv_dumper_20;
    upc_loop_monitor #(1) upc_loop_monitor_20;
    upc_loop_intf#(1) upc_loop_intf_21(clock,reset);
    assign upc_loop_intf_21.cur_state = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_VITIS_LOOP_420_10_fu_1009.ap_CS_fsm;
    assign upc_loop_intf_21.iter_start_state = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_VITIS_LOOP_420_10_fu_1009.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_21.iter_end_state = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_VITIS_LOOP_420_10_fu_1009.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_21.quit_state = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_VITIS_LOOP_420_10_fu_1009.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_21.iter_start_block = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_VITIS_LOOP_420_10_fu_1009.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_21.iter_end_block = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_VITIS_LOOP_420_10_fu_1009.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_21.quit_block = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_VITIS_LOOP_420_10_fu_1009.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_21.iter_start_enable = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_VITIS_LOOP_420_10_fu_1009.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_21.iter_end_enable = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_VITIS_LOOP_420_10_fu_1009.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_21.quit_enable = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_VITIS_LOOP_420_10_fu_1009.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_21.loop_start = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_VITIS_LOOP_420_10_fu_1009.ap_start;
    assign upc_loop_intf_21.loop_ready = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_VITIS_LOOP_420_10_fu_1009.ap_ready;
    assign upc_loop_intf_21.loop_done = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_VITIS_LOOP_420_10_fu_1009.ap_done_int;
    assign upc_loop_intf_21.loop_continue = 1'b1;
    assign upc_loop_intf_21.quit_at_end = 1'b0;
    assign upc_loop_intf_21.finish = finish;
    csv_file_dump upc_loop_csv_dumper_21;
    upc_loop_monitor #(1) upc_loop_monitor_21;
    upc_loop_intf#(1) upc_loop_intf_22(clock,reset);
    assign upc_loop_intf_22.cur_state = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_VITIS_LOOP_373_5_fu_1016.ap_CS_fsm;
    assign upc_loop_intf_22.iter_start_state = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_VITIS_LOOP_373_5_fu_1016.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_22.iter_end_state = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_VITIS_LOOP_373_5_fu_1016.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_22.quit_state = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_VITIS_LOOP_373_5_fu_1016.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_22.iter_start_block = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_VITIS_LOOP_373_5_fu_1016.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_22.iter_end_block = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_VITIS_LOOP_373_5_fu_1016.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_22.quit_block = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_VITIS_LOOP_373_5_fu_1016.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_22.iter_start_enable = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_VITIS_LOOP_373_5_fu_1016.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_22.iter_end_enable = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_VITIS_LOOP_373_5_fu_1016.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_22.quit_enable = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_VITIS_LOOP_373_5_fu_1016.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_22.loop_start = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_VITIS_LOOP_373_5_fu_1016.ap_start;
    assign upc_loop_intf_22.loop_ready = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_VITIS_LOOP_373_5_fu_1016.ap_ready;
    assign upc_loop_intf_22.loop_done = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_VITIS_LOOP_373_5_fu_1016.ap_done_int;
    assign upc_loop_intf_22.loop_continue = 1'b1;
    assign upc_loop_intf_22.quit_at_end = 1'b0;
    assign upc_loop_intf_22.finish = finish;
    csv_file_dump upc_loop_csv_dumper_22;
    upc_loop_monitor #(1) upc_loop_monitor_22;
    upc_loop_intf#(1) upc_loop_intf_23(clock,reset);
    assign upc_loop_intf_23.cur_state = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_VITIS_LOOP_391_6_VITIS_LOOP_392_7_fu_1058.ap_CS_fsm;
    assign upc_loop_intf_23.iter_start_state = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_VITIS_LOOP_391_6_VITIS_LOOP_392_7_fu_1058.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_23.iter_end_state = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_VITIS_LOOP_391_6_VITIS_LOOP_392_7_fu_1058.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_23.quit_state = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_VITIS_LOOP_391_6_VITIS_LOOP_392_7_fu_1058.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_23.iter_start_block = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_VITIS_LOOP_391_6_VITIS_LOOP_392_7_fu_1058.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_23.iter_end_block = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_VITIS_LOOP_391_6_VITIS_LOOP_392_7_fu_1058.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_23.quit_block = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_VITIS_LOOP_391_6_VITIS_LOOP_392_7_fu_1058.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_23.iter_start_enable = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_VITIS_LOOP_391_6_VITIS_LOOP_392_7_fu_1058.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_23.iter_end_enable = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_VITIS_LOOP_391_6_VITIS_LOOP_392_7_fu_1058.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_23.quit_enable = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_VITIS_LOOP_391_6_VITIS_LOOP_392_7_fu_1058.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_23.loop_start = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_VITIS_LOOP_391_6_VITIS_LOOP_392_7_fu_1058.ap_start;
    assign upc_loop_intf_23.loop_ready = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_VITIS_LOOP_391_6_VITIS_LOOP_392_7_fu_1058.ap_ready;
    assign upc_loop_intf_23.loop_done = AESL_inst_TOP.grp_KBEST_fu_461.grp_KBEST_Pipeline_VITIS_LOOP_391_6_VITIS_LOOP_392_7_fu_1058.ap_done_int;
    assign upc_loop_intf_23.loop_continue = 1'b1;
    assign upc_loop_intf_23.quit_at_end = 1'b1;
    assign upc_loop_intf_23.finish = finish;
    csv_file_dump upc_loop_csv_dumper_23;
    upc_loop_monitor #(1) upc_loop_monitor_23;

    sample_manager sample_manager_inst;

initial begin
    sample_manager_inst = new;



    mstatus_csv_dumper_1 = new("./module_status1.csv");
    module_monitor_1 = new(module_intf_1,mstatus_csv_dumper_1);
    mstatus_csv_dumper_2 = new("./module_status2.csv");
    module_monitor_2 = new(module_intf_2,mstatus_csv_dumper_2);
    mstatus_csv_dumper_3 = new("./module_status3.csv");
    module_monitor_3 = new(module_intf_3,mstatus_csv_dumper_3);
    mstatus_csv_dumper_4 = new("./module_status4.csv");
    module_monitor_4 = new(module_intf_4,mstatus_csv_dumper_4);
    mstatus_csv_dumper_5 = new("./module_status5.csv");
    module_monitor_5 = new(module_intf_5,mstatus_csv_dumper_5);
    mstatus_csv_dumper_6 = new("./module_status6.csv");
    module_monitor_6 = new(module_intf_6,mstatus_csv_dumper_6);
    mstatus_csv_dumper_7 = new("./module_status7.csv");
    module_monitor_7 = new(module_intf_7,mstatus_csv_dumper_7);
    mstatus_csv_dumper_8 = new("./module_status8.csv");
    module_monitor_8 = new(module_intf_8,mstatus_csv_dumper_8);
    mstatus_csv_dumper_9 = new("./module_status9.csv");
    module_monitor_9 = new(module_intf_9,mstatus_csv_dumper_9);
    mstatus_csv_dumper_10 = new("./module_status10.csv");
    module_monitor_10 = new(module_intf_10,mstatus_csv_dumper_10);
    mstatus_csv_dumper_11 = new("./module_status11.csv");
    module_monitor_11 = new(module_intf_11,mstatus_csv_dumper_11);
    mstatus_csv_dumper_12 = new("./module_status12.csv");
    module_monitor_12 = new(module_intf_12,mstatus_csv_dumper_12);
    mstatus_csv_dumper_13 = new("./module_status13.csv");
    module_monitor_13 = new(module_intf_13,mstatus_csv_dumper_13);
    mstatus_csv_dumper_14 = new("./module_status14.csv");
    module_monitor_14 = new(module_intf_14,mstatus_csv_dumper_14);
    mstatus_csv_dumper_15 = new("./module_status15.csv");
    module_monitor_15 = new(module_intf_15,mstatus_csv_dumper_15);
    mstatus_csv_dumper_16 = new("./module_status16.csv");
    module_monitor_16 = new(module_intf_16,mstatus_csv_dumper_16);
    mstatus_csv_dumper_17 = new("./module_status17.csv");
    module_monitor_17 = new(module_intf_17,mstatus_csv_dumper_17);
    mstatus_csv_dumper_18 = new("./module_status18.csv");
    module_monitor_18 = new(module_intf_18,mstatus_csv_dumper_18);
    mstatus_csv_dumper_19 = new("./module_status19.csv");
    module_monitor_19 = new(module_intf_19,mstatus_csv_dumper_19);
    mstatus_csv_dumper_20 = new("./module_status20.csv");
    module_monitor_20 = new(module_intf_20,mstatus_csv_dumper_20);
    mstatus_csv_dumper_21 = new("./module_status21.csv");
    module_monitor_21 = new(module_intf_21,mstatus_csv_dumper_21);
    mstatus_csv_dumper_22 = new("./module_status22.csv");
    module_monitor_22 = new(module_intf_22,mstatus_csv_dumper_22);
    mstatus_csv_dumper_23 = new("./module_status23.csv");
    module_monitor_23 = new(module_intf_23,mstatus_csv_dumper_23);
    mstatus_csv_dumper_24 = new("./module_status24.csv");
    module_monitor_24 = new(module_intf_24,mstatus_csv_dumper_24);
    mstatus_csv_dumper_25 = new("./module_status25.csv");
    module_monitor_25 = new(module_intf_25,mstatus_csv_dumper_25);
    mstatus_csv_dumper_26 = new("./module_status26.csv");
    module_monitor_26 = new(module_intf_26,mstatus_csv_dumper_26);
    mstatus_csv_dumper_27 = new("./module_status27.csv");
    module_monitor_27 = new(module_intf_27,mstatus_csv_dumper_27);
    mstatus_csv_dumper_28 = new("./module_status28.csv");
    module_monitor_28 = new(module_intf_28,mstatus_csv_dumper_28);
    mstatus_csv_dumper_29 = new("./module_status29.csv");
    module_monitor_29 = new(module_intf_29,mstatus_csv_dumper_29);
    mstatus_csv_dumper_30 = new("./module_status30.csv");
    module_monitor_30 = new(module_intf_30,mstatus_csv_dumper_30);
    mstatus_csv_dumper_31 = new("./module_status31.csv");
    module_monitor_31 = new(module_intf_31,mstatus_csv_dumper_31);
    mstatus_csv_dumper_32 = new("./module_status32.csv");
    module_monitor_32 = new(module_intf_32,mstatus_csv_dumper_32);
    mstatus_csv_dumper_33 = new("./module_status33.csv");
    module_monitor_33 = new(module_intf_33,mstatus_csv_dumper_33);
    mstatus_csv_dumper_34 = new("./module_status34.csv");
    module_monitor_34 = new(module_intf_34,mstatus_csv_dumper_34);
    mstatus_csv_dumper_35 = new("./module_status35.csv");
    module_monitor_35 = new(module_intf_35,mstatus_csv_dumper_35);
    mstatus_csv_dumper_36 = new("./module_status36.csv");
    module_monitor_36 = new(module_intf_36,mstatus_csv_dumper_36);
    mstatus_csv_dumper_37 = new("./module_status37.csv");
    module_monitor_37 = new(module_intf_37,mstatus_csv_dumper_37);
    mstatus_csv_dumper_38 = new("./module_status38.csv");
    module_monitor_38 = new(module_intf_38,mstatus_csv_dumper_38);
    mstatus_csv_dumper_39 = new("./module_status39.csv");
    module_monitor_39 = new(module_intf_39,mstatus_csv_dumper_39);
    mstatus_csv_dumper_40 = new("./module_status40.csv");
    module_monitor_40 = new(module_intf_40,mstatus_csv_dumper_40);
    mstatus_csv_dumper_41 = new("./module_status41.csv");
    module_monitor_41 = new(module_intf_41,mstatus_csv_dumper_41);
    mstatus_csv_dumper_42 = new("./module_status42.csv");
    module_monitor_42 = new(module_intf_42,mstatus_csv_dumper_42);

    pp_loop_csv_dumper_1 = new("./pp_loop_status1.csv");
    pp_loop_monitor_1 = new(pp_loop_intf_1,pp_loop_csv_dumper_1);


    seq_loop_csv_dumper_1 = new("./seq_loop_status1.csv");
    seq_loop_monitor_1 = new(seq_loop_intf_1,seq_loop_csv_dumper_1);
    seq_loop_csv_dumper_2 = new("./seq_loop_status2.csv");
    seq_loop_monitor_2 = new(seq_loop_intf_2,seq_loop_csv_dumper_2);
    seq_loop_csv_dumper_3 = new("./seq_loop_status3.csv");
    seq_loop_monitor_3 = new(seq_loop_intf_3,seq_loop_csv_dumper_3);
    seq_loop_csv_dumper_4 = new("./seq_loop_status4.csv");
    seq_loop_monitor_4 = new(seq_loop_intf_4,seq_loop_csv_dumper_4);
    seq_loop_csv_dumper_5 = new("./seq_loop_status5.csv");
    seq_loop_monitor_5 = new(seq_loop_intf_5,seq_loop_csv_dumper_5);
    seq_loop_csv_dumper_6 = new("./seq_loop_status6.csv");
    seq_loop_monitor_6 = new(seq_loop_intf_6,seq_loop_csv_dumper_6);
    seq_loop_csv_dumper_7 = new("./seq_loop_status7.csv");
    seq_loop_monitor_7 = new(seq_loop_intf_7,seq_loop_csv_dumper_7);
    seq_loop_csv_dumper_8 = new("./seq_loop_status8.csv");
    seq_loop_monitor_8 = new(seq_loop_intf_8,seq_loop_csv_dumper_8);
    seq_loop_csv_dumper_9 = new("./seq_loop_status9.csv");
    seq_loop_monitor_9 = new(seq_loop_intf_9,seq_loop_csv_dumper_9);
    seq_loop_csv_dumper_10 = new("./seq_loop_status10.csv");
    seq_loop_monitor_10 = new(seq_loop_intf_10,seq_loop_csv_dumper_10);
    seq_loop_csv_dumper_11 = new("./seq_loop_status11.csv");
    seq_loop_monitor_11 = new(seq_loop_intf_11,seq_loop_csv_dumper_11);
    seq_loop_csv_dumper_12 = new("./seq_loop_status12.csv");
    seq_loop_monitor_12 = new(seq_loop_intf_12,seq_loop_csv_dumper_12);
    seq_loop_csv_dumper_13 = new("./seq_loop_status13.csv");
    seq_loop_monitor_13 = new(seq_loop_intf_13,seq_loop_csv_dumper_13);
    seq_loop_csv_dumper_14 = new("./seq_loop_status14.csv");
    seq_loop_monitor_14 = new(seq_loop_intf_14,seq_loop_csv_dumper_14);

    upc_loop_csv_dumper_1 = new("./upc_loop_status1.csv");
    upc_loop_monitor_1 = new(upc_loop_intf_1,upc_loop_csv_dumper_1);
    upc_loop_csv_dumper_2 = new("./upc_loop_status2.csv");
    upc_loop_monitor_2 = new(upc_loop_intf_2,upc_loop_csv_dumper_2);
    upc_loop_csv_dumper_3 = new("./upc_loop_status3.csv");
    upc_loop_monitor_3 = new(upc_loop_intf_3,upc_loop_csv_dumper_3);
    upc_loop_csv_dumper_4 = new("./upc_loop_status4.csv");
    upc_loop_monitor_4 = new(upc_loop_intf_4,upc_loop_csv_dumper_4);
    upc_loop_csv_dumper_5 = new("./upc_loop_status5.csv");
    upc_loop_monitor_5 = new(upc_loop_intf_5,upc_loop_csv_dumper_5);
    upc_loop_csv_dumper_6 = new("./upc_loop_status6.csv");
    upc_loop_monitor_6 = new(upc_loop_intf_6,upc_loop_csv_dumper_6);
    upc_loop_csv_dumper_7 = new("./upc_loop_status7.csv");
    upc_loop_monitor_7 = new(upc_loop_intf_7,upc_loop_csv_dumper_7);
    upc_loop_csv_dumper_8 = new("./upc_loop_status8.csv");
    upc_loop_monitor_8 = new(upc_loop_intf_8,upc_loop_csv_dumper_8);
    upc_loop_csv_dumper_9 = new("./upc_loop_status9.csv");
    upc_loop_monitor_9 = new(upc_loop_intf_9,upc_loop_csv_dumper_9);
    upc_loop_csv_dumper_10 = new("./upc_loop_status10.csv");
    upc_loop_monitor_10 = new(upc_loop_intf_10,upc_loop_csv_dumper_10);
    upc_loop_csv_dumper_11 = new("./upc_loop_status11.csv");
    upc_loop_monitor_11 = new(upc_loop_intf_11,upc_loop_csv_dumper_11);
    upc_loop_csv_dumper_12 = new("./upc_loop_status12.csv");
    upc_loop_monitor_12 = new(upc_loop_intf_12,upc_loop_csv_dumper_12);
    upc_loop_csv_dumper_13 = new("./upc_loop_status13.csv");
    upc_loop_monitor_13 = new(upc_loop_intf_13,upc_loop_csv_dumper_13);
    upc_loop_csv_dumper_14 = new("./upc_loop_status14.csv");
    upc_loop_monitor_14 = new(upc_loop_intf_14,upc_loop_csv_dumper_14);
    upc_loop_csv_dumper_15 = new("./upc_loop_status15.csv");
    upc_loop_monitor_15 = new(upc_loop_intf_15,upc_loop_csv_dumper_15);
    upc_loop_csv_dumper_16 = new("./upc_loop_status16.csv");
    upc_loop_monitor_16 = new(upc_loop_intf_16,upc_loop_csv_dumper_16);
    upc_loop_csv_dumper_17 = new("./upc_loop_status17.csv");
    upc_loop_monitor_17 = new(upc_loop_intf_17,upc_loop_csv_dumper_17);
    upc_loop_csv_dumper_18 = new("./upc_loop_status18.csv");
    upc_loop_monitor_18 = new(upc_loop_intf_18,upc_loop_csv_dumper_18);
    upc_loop_csv_dumper_19 = new("./upc_loop_status19.csv");
    upc_loop_monitor_19 = new(upc_loop_intf_19,upc_loop_csv_dumper_19);
    upc_loop_csv_dumper_20 = new("./upc_loop_status20.csv");
    upc_loop_monitor_20 = new(upc_loop_intf_20,upc_loop_csv_dumper_20);
    upc_loop_csv_dumper_21 = new("./upc_loop_status21.csv");
    upc_loop_monitor_21 = new(upc_loop_intf_21,upc_loop_csv_dumper_21);
    upc_loop_csv_dumper_22 = new("./upc_loop_status22.csv");
    upc_loop_monitor_22 = new(upc_loop_intf_22,upc_loop_csv_dumper_22);
    upc_loop_csv_dumper_23 = new("./upc_loop_status23.csv");
    upc_loop_monitor_23 = new(upc_loop_intf_23,upc_loop_csv_dumper_23);

    sample_manager_inst.add_one_monitor(module_monitor_1);
    sample_manager_inst.add_one_monitor(module_monitor_2);
    sample_manager_inst.add_one_monitor(module_monitor_3);
    sample_manager_inst.add_one_monitor(module_monitor_4);
    sample_manager_inst.add_one_monitor(module_monitor_5);
    sample_manager_inst.add_one_monitor(module_monitor_6);
    sample_manager_inst.add_one_monitor(module_monitor_7);
    sample_manager_inst.add_one_monitor(module_monitor_8);
    sample_manager_inst.add_one_monitor(module_monitor_9);
    sample_manager_inst.add_one_monitor(module_monitor_10);
    sample_manager_inst.add_one_monitor(module_monitor_11);
    sample_manager_inst.add_one_monitor(module_monitor_12);
    sample_manager_inst.add_one_monitor(module_monitor_13);
    sample_manager_inst.add_one_monitor(module_monitor_14);
    sample_manager_inst.add_one_monitor(module_monitor_15);
    sample_manager_inst.add_one_monitor(module_monitor_16);
    sample_manager_inst.add_one_monitor(module_monitor_17);
    sample_manager_inst.add_one_monitor(module_monitor_18);
    sample_manager_inst.add_one_monitor(module_monitor_19);
    sample_manager_inst.add_one_monitor(module_monitor_20);
    sample_manager_inst.add_one_monitor(module_monitor_21);
    sample_manager_inst.add_one_monitor(module_monitor_22);
    sample_manager_inst.add_one_monitor(module_monitor_23);
    sample_manager_inst.add_one_monitor(module_monitor_24);
    sample_manager_inst.add_one_monitor(module_monitor_25);
    sample_manager_inst.add_one_monitor(module_monitor_26);
    sample_manager_inst.add_one_monitor(module_monitor_27);
    sample_manager_inst.add_one_monitor(module_monitor_28);
    sample_manager_inst.add_one_monitor(module_monitor_29);
    sample_manager_inst.add_one_monitor(module_monitor_30);
    sample_manager_inst.add_one_monitor(module_monitor_31);
    sample_manager_inst.add_one_monitor(module_monitor_32);
    sample_manager_inst.add_one_monitor(module_monitor_33);
    sample_manager_inst.add_one_monitor(module_monitor_34);
    sample_manager_inst.add_one_monitor(module_monitor_35);
    sample_manager_inst.add_one_monitor(module_monitor_36);
    sample_manager_inst.add_one_monitor(module_monitor_37);
    sample_manager_inst.add_one_monitor(module_monitor_38);
    sample_manager_inst.add_one_monitor(module_monitor_39);
    sample_manager_inst.add_one_monitor(module_monitor_40);
    sample_manager_inst.add_one_monitor(module_monitor_41);
    sample_manager_inst.add_one_monitor(module_monitor_42);
    sample_manager_inst.add_one_monitor(pp_loop_monitor_1);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_1);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_2);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_3);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_4);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_5);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_6);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_7);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_8);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_9);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_10);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_11);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_12);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_13);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_14);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_1);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_2);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_3);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_4);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_5);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_6);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_7);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_8);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_9);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_10);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_11);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_12);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_13);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_14);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_15);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_16);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_17);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_18);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_19);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_20);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_21);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_22);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_23);
    
    fork
        sample_manager_inst.start_monitor();
        last_transaction_done;
    join
    disable fork;

    sample_manager_inst.start_dump();
end

    task last_transaction_done();
        wait(reset == 0);
        while(1) begin
            if (finish == 1'b1)
                break;
            else
                @(posedge clock);
        end
    endtask


endmodule
